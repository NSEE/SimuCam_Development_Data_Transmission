// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:48 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BptTANKd4bHdLqC7xR1S8R1BpGHXbCfx4Ub/U2nrGvB0p6pS4KCeJlUk0KqjR9qQ
p7pOb/P/DGDYSKdW6uUSwBJPuPl94+qkNz5ARCJF0WQqCIoqbB6u0irct+e5BuRW
vye7+JK11z23xdjNnTvLUEfCapNuYImXeuBiv69h428=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5728)
WBwJ/CguiDl6UnjvbMeKDwX0n+lR7Dth1YjlorcQpJiXZnBWU4652VqYCgO436SY
8LjwWdqyV8CozIo/ZHac+zNf2Z2Tcx4IXf9bw3pg+vUftWqPfNiMwk0wOrF0MYyc
wcDPoCw0o+qhrTQ2xzgq/EAGzgZbwWCvHpiybzrFMUF24mJt2UdoEJu0q+a/bvSo
Hd4OHFfH7yuNVPQmc5jO6uRMqO7F9LE21mCBIz1Nw57XhJR3nQQs/KG6oNlrM/wY
8+mNNSJFuYnBcSlJWWzdU1ioKkF0yWVLp17zOpvWHJw6AMa6TLR4m40dMDbicJ6z
8DXjds3E+2uw9i3zXOT97/iJkYJmbpVs1jC+ivtWK951bZT3VYrGtKxZuY16ODhH
kvmz/baCZaqhywMQImYrx/FWSDl5baqZCyBNdlhM99Ka9wfX4eSfVssbOomTsMH0
R266n3pWgMIwLoXCHmoEuhULS5R4wmOWpAV1mad9HeNaGMrlZ25j6sioryUpkdxf
9h7DtCrDibur+ZREv05d5pGkSHKFnHHVxrZ0jLGP/FPUdVo4fMVnn+SPq6XOjA4E
1RnRE+SDIHeAc6D0Kfj+xEVJRbGQLnZPDhj6Qraa6gaQKWybXtC5XgrDDxBmvK64
d1TDjpk/lo3VpRyod52CKu8QTy55D/pUOvAyE4gL2/+GnHk8gk8gncbHpC0YOk7u
547Zug91uuJSKKIMJ2XXk09tBy/BNWXmWW6WMjAM+LxxWlseXojLzDD2fOd2DsQ9
W6zGoT9XLrW0ZmJYOf0Ir0g23rFLvrMyBEhfqiKoSmxjSnptJA2ROEaonDs8cOUL
mDUJGqPiJxtFJXpQHHNf/K12z3B8tkCwnXOlMHh00Yg+KqyHc36jYOAahuk4g8+W
WU6NEwwqddaOy+poYTmFj8hQUFhExrS2N5+Z/MuubgMZQBZhqdvXmQxdV+3JUlYa
hHBiP40WjdtbI2d08SyfGlZHTkE7N/FEQu1Na4GhOGu6WMDHoQDGB679APhcL6LA
NZ4L5XscpBE8d44lSnsurDTyD/Gpd01y99QAK6JcZ2wgC4ZMelanR39gQm96sGQj
epFx8TARmclZjeq6AfxqG5WgDoLgdS+sOCILcgrxN/qhVdQL1MkqL18TOyI/wYHH
SvkjxjhUG6benflP6eB17QMYOF+2OxUjvt7Koumpv6MSo2gVbC0u2mmVecBPJnJ/
rWwCwmVygyKmM+nTCMZFe003eWNdfG32zucgOcA5o81Gp2PzsW2R2k5rpQ1TrxGv
d0HuYCEjb+x7H8hcQ+XAmLjck9Go36m6u43ZAGxqx9sHn7n+XKDxAmQ+1WykMGBP
cTp/CQcl5+EXsW550c3XRRbaOBqnlIH3mlYRX36/T6h1CcGs+fry3d6pfh/82bsQ
5tAWuYyLH24RqGf5GFqQYA8DUce9Mj/EpHOO9x2lfiso6OiUhIpJeqhpBJZTdlG8
LddlaIPpJGFgmaJjrePaMdOkx5xgyIOryu3wY66j2MTp6DNMsWbsM5LQXZ4Y+POG
G0vM2iamSqtVEWoGetKaxZ+X3Cd9/a1rpLLahRytFaAzyUTWdNFZXoNnQvCf8wE7
fZ5sqEeIANFgZl+e94MR91EFhZrOMuG0LT4zJ0b+FSYaG5kOuxk/1lpeUgSM7VFB
drLdPvlM15rIwDE2I3vHar6pMS2Kzfe2tipIIcQW5NvQPUd/15K5UCG/fA+Op8iZ
LWPVlGGal/6Soi9KxwU2hulzcHE1mhk495VibU07l9JwOLTVULag5H6GR4D2fmLt
1FaswmSngaemTdyFGCXFcXRqOfHJcYDlj4IgttZXk1keBEVduD1VB2aOq8vpSSCK
6XNWflvD6akpaiONyYLFvPchrGOC1hPpF8TRvxHspxuXWCq4V3FECOElhpP8atxG
Z3suhc8msLYyCqbk63ZknJB4nBOS8kgI9XBD7uk5Q+1JvCUijJ6tBX+O8G/ChM4S
tXRA4CbmTPl57iHLxcaQiBkKrWFPpRH23aQBVFgYSNUoM2xuofRb3GI13vvVBu0E
nSgKy9OyowllKjEJ5pqvFODHnlxjLLFWxR0T3grBMpspjp7ILSDPsmbihCIjRj/X
pC13HMSDONI58Qhtgkwjn7x5shE8fnyzf3zosrK5MjSVdrDtpZThZK+PcK6IrGOu
4c8ku5C061GdbkGpcLLW4dL9RKw2dlfoVEsMY3dAL/x/+fffqfZu9BjYK8BTKueT
Wm0NJTcX8s3HAol1Vnz9rW4IB+CaIwWeBeV6V5GfbG6chqYbB9T+aJaBtH53VLlW
CsWUsI/uXZEqAIfj6fTbUbTLeF/DOCjcPyu7nwM/1TF3sil3OKBELXyPWEbExO2d
MVNS9zcFm5VsEPjlutH4NdS8ZEwJok3cJaQvRXFauhf2Fg/T+xGSGno73ariPbXj
VwKQpIWCz8jfKys7hfPuut6ggGeqUdlME2JhoSutOPs1/7PatlhMYD6XYuYsIIev
6Kaw3fucrqpK1Z1tPQSukH6DsP8XsFO4EFZBaDD47LQ5EDWGDHFhmFv+TTibcYem
cLI+K9o5/6T+kUrC1a1WtuBIDH7pAoA1LHTh1uv5pEdG8ZxGdN1rNF75qmpBtmc3
09z8pK1m7chjR99nlmXOVhKh+0g/0t2DgQww3fy74TgzEqtE2HZQK3qWhhvwLrd5
hNu8B/8TmxzIaOqBs0+hx6zJxbUb+2bdMYnamSLrtSNhjfffLzH5DhMJFzz0tXF1
D7zfGtW8X7Lhs8OJolsmTMAMebb8W94WxKhuyn0I5RGu5trpafs5AkXHZCnET1dG
oyFb5XrEo8GthfEpOe9zQ/5ry1yLiTXfR8u9RWU7oSS5rEKpKkN8KPptXe7cDHCj
3fCI1Ta/b1ZjsUbAibxYXeVExH4e3u+/16sPY1AuaUS1eHnIzpprAfwOCfRxedBy
/4Gt/y/pjPgiEyJqpPu9WypGdviw1GiiJbbk8mOo3nQKXLbTpgORIEXMXgN4elke
v9jEZCredwk2KnNu6rdfP3uhP3ZP6FANEfwA5NNGfv/Z0lbn/AMQXHbLTFlYlJVJ
dotlOukrKt+LhQvc5gCtXUmlYrcrvyMJfQRQh/BkNFByo2YAlqBpeS2i0nm7rHqg
j/s3ImhCTwytC8YKcka4duhoUV/PevYXtM88Y/JMzGwXFHmwdiAD4Mr2l7cXqYOi
MjuVAz4gWDyehN5gWp+DfdZia2xiPZIn319DX02OBg7Drs4mCRImy5Jp0QlANoSr
vlV2eu2WldUSzLvA67AOFpeKG/o056hS84jXlp5Om4G5S8aR8udYaELd2mWl9tPz
yYCiNZHxC1AIkba4/OJOWn4StBnPIsW16Y103mwUP5YCvqgpRHzQzHzB0rdi6kzo
0HmDQ3YiBZjLukDLC4J83vvVT4G4Op914gzRq1TUcybIkTQvXDrqzdhQlVXiNRWV
/rqHs0TEJqUkAmltGq4EP5APit0No0h4hFndwk+m0Ugqgk46lm9V4HcR20Fc8VuF
968SA6ehjVRkGvSAOaK2o4+epeR8hts6SaEmzaYIHQOgrOMDtkQE8UTtL1vFp29P
qhQLyqd2JEK+z886T7BVaHDjcaTOKiMu5kQdqDOWPLmSVJeQBNs7d/Mw0yodTBje
i4hcF9R2KaGL7+QReZpjeixMAyAgZRvsEp0hat3q23/UR992EjIoiHtW6HW4J3Sl
ZtvkCsqmiZ4ouESpTs/n5ijhQOc2/NY+4JK2P0t8XF3Bo9UqM3ErIW8p345OvJfD
OIQ4d4SLSfGqxbwRWzMnYMbRmNqyw5HfvozlJQQp5hTi4WyRDKvQ0pQ6kXuJIOgC
w6F0fHO8ci9swIyk4BQ2r0oJJm0QJ41iSCJoKQDgEdbnRTaPe/YXkiKIKPvwe2Af
5uQWv2WYiXfVenRiwAA374O8eVPKL9xgSvF8kdAbEtXbrzBjGAEbCphJc8xx6pvI
2vl9/qU33aMBYBtZaMNzclJBPUDAu76iLs2SRTRpCP8gGgTaSZrSyNHGjH4wyA5j
ytN1ERpngWOfl8FHal21g+HgrQiYOjAbku2CKeB+aIzYVM9ugCJjdy4k/zPgNUfo
prJ2HdBOrmDD/lAHHXpJahLEzUuIK/9mxDsavg6s5p7Oqm05Yx33iv8ey3EYD3JW
rfeeFNdcrCtsS/hhW7ZJ/DXlDdde9GhE6+yQDMxapj/Z+FIArWuE33HvBxtgzacW
in0okB3EAvIwThluorL4dPFiPkS7Ez/y6w7C6fIIcH7ufBUbBbDdePVkPPA6Y/vZ
/eT8dUFxmxmBGs/TpRgbzQyLv3z2436BEbSS3pYq1ES5ZTM1SfiBb6H1umyHE8cv
HsRMvySmkbHE3sPg7oe2mMdslcWf4MM/I6vBxbxh27I8C/Sxuw6bIx46nWvWaQpY
vewO28iL1xWimDKfpV1g3p+DoY0U7y0YQ48x7p3BdA+P8l/j0lVblBD4/JxISPTI
xgKt3fen9wxAlxf6B6fC0MNLepw3GuecqqjWsgNoxdT7o4F+E7Bun8IkZD21wkKU
cTlZtsPZhu9cN60SCxCZZc7VPUcNoauhnS1P88yY7Mo7T1e0VbpnqKDSXOYGKPpF
v37oqrzn+S22eux2pn8AuH2aqBtHuZXqTnSZDTGjeyLa5nfkB7pWaV7xesjDaPQS
ec5tCZUaldL06xF2n+g33SPgsMoeo24eUYnW8Po6XDrPBK2amr/75v4X1ByT0rYO
kMBDX1HLUwg3/dFp4mEbrizNGUB2lj/FtbEPHg/opk2D/o1TF79xxiwHnn7ryeKp
QSh4YlLGtds/jCu1G//1yPIz2GOPyc/8UN53QQEIegniS1lYhxzWlWzmHdlazPkq
P5eeRcA6xNuW+cBz0C4TflR+8TSqQfvAc4H4Am57oiWR0NpOzDZaDVgRfhAqjKPD
zv1YKgbfS4JbTQAAFxS2btL4oaqxdesNtKm01f2ADMjLJuqnpP3vCOTckB3xpF7D
6OI6VLa6a+UxEn3RxDjnAeSCREtThnYTrvFowE7fkv58fv6W+gZLDzBjBSLQC/13
vfL93Nbg9YnPQTkZQjvF8DLMz41SzCc+a2ItAWRbD0Gufu/Ke/MQjOjPANQt/JNc
MXcBwhlHA8OMRrgRb4GeAq6zm1y+4yJtqNhF1/Wf4UX3EHAnuoUC8cLeFNIReRXS
/ugVfN90KshMYE2NbrELywWHk+31PvkwiJaJ3ahjD0j1X4saAbHBXEa3C1V5vqPV
6UYjV2HdOAqp/WlvdVsp4tsRrgw8Nabl5YTa4aJOD/Cg691rYzHdf7WYnJm9TXGn
KVxG0ky5IZ6WDT7H7Kc3iVAyOeH344RLogAdm7FTy0cooKpWEpFHtR/rkLdlopne
mHmcTa4oFoXTqlZg7CCtVGRxs3cuCA5TMU/SBZd52oUjs1SwSrBelK3JHRpM6HH3
S0o0Jt/Nfr8Sg+DRWHv4teLY160t5VJkZFnSAjnzzpIZP6LkjPxsuiPQ8RxWwt7p
qSaWgNh9qWWbKX6arCYbT53gG/JPnHPgECclP+gAx2QQ5PI9bisOnlcb2stzZbUb
ZHOTHjir05KpxpdEUBCCHrzDfZUge8Ogdy5urNjBbqm5undB15MROamSBEqhfCqP
t0AroXl4jjBw9JxOnZX/6xGn5QUHXhIbZ3B3PfQiUjr5Aq3E0+J9ieTTTXkmpe2a
nL96ANYdQqsJgCJT3lTNqKPkZ0b1lJBISfr1puCFTBvl8UzF23PNaZ9y1mYukaax
BMtnZLNqBAtma4R128uaTlGfEkSHiVxhuDLVhUvriGDb4QAHjHSr5PdErRK3TxoM
qAbgEcRAh7uDU55A1SzSU6yW2XB4SjzayIWl4fzOaY3Ome+RI8XTJknxT9u4wyAK
ZZrDdv/yzsyVSpQ8fl4Nki707uBuxsM9HP0w95zGjuOGgXV8NQdREKm7wqZbB+1E
l/LKMdVbhrHgx/H9yVWExUj4FA9SswGUcmWWoghH8rg9bl1gGzI06sGIVdKuerDg
+TzmX4woej7k4OXEPMr3i603lCFMemelNzF+kf74N5dg7uwWMUiGzD4hF04ITCpJ
2+NPQlZK4i0hhqe3i18SwGpGjLx+iiDQOSSRyOO400DX3i2gxFeT6Sb3Gj2fTefp
vkoLilKwf9rW/DMR4D1okTz6jddgTrqozblx0wnYa9N41dDXVrNofQdFdR/esDYp
sw7in7IgaHvTft4KDRut1Ls6sJ/yN2RJLc4nGbyB7GFwgXHeLcbevavYKJjSj3iP
35AS23vjVx1BOrbyXAQVk6JivcZJk/baHxmTYNv3kTuifuCASS/txXXhFdqyPFnl
jDOLWqheHpuN5RxGIOsRzNDrHQXmXP4Kjzg51eIyrC4onCLbM820trhPI2j0SN9v
Bs09RXQItCpxjuuPiXuRdhdlK4YTwjvahii/fjgRq5kZ9616gw57XajeVgaiFc6A
XcXXqQtNdyKUS/RrM4qPYlYRdroBFfqhT9YtZHQVJelSxPmLny09XHX12a7lvjst
DIVDHa5ZbmdwI7wonilVEQ72Uu2Vnj+OlhotTCtZ07OEUzDUuLAq/pubQ1uZQ2P7
Q+q06filmtxrVEIp2L1+W4nvju4pGyIXoPIDdXwx++N1q2PKSUNLnJDbbmUEeXKd
mZIe+BbOhfboYbKSM42Jkktwq174qu7P/BD4R/pbWPVGTPkCTbGjJD4duaVv2XYn
hbViPw/CSPn/seTY8ImYo/xoR+voaBzIyI/4x5wYB8DYWKfgLuCw4Qa6Skkke1ji
Nn0lLD3rJi0+glh9Aw8dNe8yjjF24fydz2n+O3mWj7LjXp422CW74AgzxHPJ8H9k
gHZpcdkk45nMHzDyeFUxwM7XlkJh/uz6GPRrD+z8NTzNT9IIVCUrcTxmzAR19qH9
YoXffmGDWj+i6cJmMAiTO+YpLTvlrB9FkfGNJH2ElibB5br7kNZZwJ4QjGvbt4p0
AA7SV25iptQPmndgZD8y//JI+j+XhOX5Ml487BBvuuwJmp4Oj/COGerUhO1N8Pk0
puCYT6hQj5twyE0QuKv/76QwJB3lTTGEN0leweWNEDQOVgksaHyphnYrtACueuP0
/vCQnrDk6uSpTb6dSa1WAozs2TxKFnkyXD11qDq4tG9BYhkCFtBoXSbw0qCRr78G
MiCR3mJfZKkwGprllmNy1yRPRjXDixWXwExp5ZdcM5F3f3Cnm39bxJZBwgP9JdiL
1StpB5f89OFmbi1yKZk5zVxzNJ1eqS4kdjolF4BwdkP8V5d6SsZq3A9iaip6isgs
MAWqWyiaJj9WSmk7oBEejU3vPKa5DQUnoxZ21EcHrB7C9ahXe+BpDPvI2G1LyLEs
9hAQu1w5ASmvcA6gE7zFOPIPWXvUihbMYhQESDmdLR5fro31dRjHSp7j6uMn7K5b
bKtJREY5SFgE7tdRYnkBIBqUVQX7dupYPBDpRY4ho+ddETTataaK2d4uwtfeoTz6
OrRcqaUHe/LD9qt8mprA1yCmssXWcq7Kt7f9CI1EwMBDAbWO/vfXLmTJBqH7VwHv
fyQSQ3omP+dNu8f6gMo40BjNWEykALhcerTSMCSnEobKKwGCJtfL/OGHAy8mnffZ
s2fKC4BVKcD0qqvpJpgBDw==
`pragma protect end_protected
