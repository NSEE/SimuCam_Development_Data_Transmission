// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:48 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PXbRnYBrN8M6gryWnrxKD7lx7wSuUrtBo/WybYGLwDS2S/VEyHN48o9oc5QHzHYp
6EZQCTxewlxYB94rINdPbhvYiBwyWyCxklqXsFeg95eF0WBvJbCGk8PmDb45bRwX
6M964LIxrNwzJQ33o0ld2ASqpSdw3P8C16oOdhvZdn8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2400)
k+Fa04WxB6WDcVn7vxPVmDAd00xqS3Pj09XSngKwmT6Uu7pEjip0uxizDYQciWXl
3t8iTg1z+CBHtQfFLQDoe9VNGNWKoLwCJlCTHFCHhpxzWkyJrL+BKzyD0JU2QVcx
DPL/HcWei9ZBtoub3oZz0Nla5vBLDVX2sUVZwRA7fdhm2GKf8ArCDsrULRXhZOOh
LWzfIDLp2QRXRCkKu2aqn5smoVG07QDxQBiV5MHgKEHruOHi6oSf1tHsvanFX2Uk
hpYJCdCcMJS8vJKwFxLgY0BzRtl+IyatM7t0I3EmB8VdDzeAOHd4ZzARo1m1kQZq
kjEqXkP2ywuQC/YCo3i110f6jD4ZFcAeUMhcTqjX1fD3IB4CDxkczu8mgo9oqAJV
wiNW3leXHB8he9b6eKKA+T6zgqNtzH4Ys7zbu9x+H8QMYyk8OdQdMznM0vhD5iBL
UtoprI4QrloWBtw+NFKNk9jXkaJ1oEJh3nFfJMkmNnwqu8pSjaGUXoTWIlV4S5rH
I2zCYdHc4inlB/kxpcLrchVIjlvmjo1mleDt7VNlwqXYe3KXWLn0vB01TYlHczDI
LlPiDdPK4Mz8cZb2akz5R1ohilz+L2356V5HHtWfhZFI2mmFTK/NueSjaXghmcRZ
7RQv4ykb8SToW1So55jIdsocfq5Hc907uxeOlz5tvtpmF82II9Whb98rLtACE20q
/kQUNj+zx7o0Ud2P0/F1rs+d/Ae1coltQVx2axbcdoFPdXPLHKhFSmfYJEzf0MtI
/AoA4d6n2rRQFtDzxDg8N8Lb7PwDavQP6EuzBBmjiBj3TpXQJF16i6hivGrfDM4U
/w7+GOkToMsDTIprvVvzTA7g5G6u/Jn7HA5rJCADJbVYJ+spfhvDu1IV9pmOXL0w
P1acJWlOE0iU6UZ6rLcH7KgB152v+cKvgmPmzNVsOKIiHZ5ElD5jKUgd9iHxUFxD
x+17RZX6jy9rGM2lCw97HxuySubhaq2v7hXNCJI5RARURduIoPwsI52cNR91ifIW
wLQx0xHEEXzOfZG5GMcOr8cOPSrwR9hsLLKUYyr/N1LMTHaPTeIZAJccs5ud7aMB
5v7i4X9MT67FHBEqpYEi4axdMU0ohjayHBzu0gNHbKXp3GCmwmWi1wH/MapIrVdS
fgPtO/Gt0lIWcIV2TexBBeirr+CsIUujb5C4yaZtWfD0GWQd+FiJ+9OiLhbV1O1C
+hxhf2fDOggJffH5ni435tnLxi02fJZaAzFvub6bORb0xpXkOcpDVwjgbNJjDcsS
V3/39OdPxHfONnmsFAxnwLly2K8AQ3ayqUA9mCuEo1c1BFYWroqJx6rYhXhVUXOM
KADnXRnSmUV1wm24kzxApOCRR0cSEUFkpAMafS55FWYcLoYAFS4ofpnHaSx+Necg
z/cjB6AU2/xHlpXascR48cY+lvZjn5Zz/0NwP1K8jFlaS3gTtCWjOaw5/O36f/+g
gAWBZYeCgrta2smwZ7E/Q/QteXQygKa2LP2ZrTmju+kIK2p60gPNZYZXwI2tOZXU
Hbsx9+DkqVez4h1RatYWyd4eWj9kqdaivK4o0BppgbbV2KfMI7FY/659wFLg9QHp
zM5Ml8hqDHcSrSa9rpDn+hRFFDtDhaFtcm9MSKkozLnuVZLeGsKzV9LRSbZEupkW
SK4VbqSkpsFjqc/rn4j/VCNsntnG6DIRP/lr/9tvZervXpaR6XjJiHQG+Naxoa1i
Ze+vfubEx/Mnu7cU+4Me5KtKcTmlJgeEc5wbNL0ms6MnqtrlXUpIvIQAk9rjvQxa
i9ar/eOPNx8yILfNlf3PXVwUeO2xlClWlHA+8LtO61I7YrtXYr1a+YcqnCAM1ncl
WypszN2GC9yowPRQg7GF32cs4uXk6M3WDZDDjiHDlplca94jKj4LNXoIJo4cr0YQ
vQelDcN8ZVtozj4Eg+usiczV4m4wqwqr7iOs4fXUViT5JjuVCcWbTCY3oOqIWKfY
cHKyfnal2N6ellRapTDzFgvIkIqstv8F/LR6LQ+anA/B64dB/qo77rnCv7FsTMjR
jP479lxnAO7m+4LnN5Tj6ym0U+njzou96kyTgO5mbTFATPHAP7RXdTIv+Vtuyfk4
1syhSo8tuKyvnocW9xom/D8DOKNfFDwrDqIyN8yaNq90F4DXP7ULIHrZmNVoWEdT
qc4SNYrcyey/gJzcc5bEp/dtQ2HFvXbs4AGqxs52mMGh2ewgTMjpw++EWxS9EGhP
Rbtbf9fHzU33+gTlB1+yTC+8zEiE1xxAGqFE+XXRggsG392qqWPe/YIaQXkpBBFr
oeVo+vQXuIa8cTs6fwIDGLfqOX3uPt/1YZ0YwQ5BOSdSzSUo1cTaJ8BZigdwjcMk
bk1RTdaQQpQyBeKHDcBS6nVkMcOMZzhV/RsAjyy/sRNV2wEQvJ1K2uyylH18QtZx
cZ1wKvSL/gWppgzTKmV+QPsCU90+PRCQNn6tUjtH03m0kHtbKhP5EnoCHwrFsJzn
epXjBR307SbC4P5aO+ViANv/Fg9hGHINXKA+R/sT1Tk2N2gVbT1uQaMJNrgSZsl9
yYcQyA24Aj/jsZ80jBDptw6+SaMJEjMTFqAhFWR+GhL0/YDrFc0luw4yNJ3uIUrf
roCbAJvT1Z035dalqFCG/D2SjqVkua6KB6Yp0RGpGBDaxtXnyRTAWFRAaS5YiHhI
NRhT8atTbz29bmEvn4qibeNWS97CWVft1CfeEKk6jCFpTnKnycRAnGi2VSjc0cKc
I3ZbHTevSvlgWElzBrK4IFk5sZVrnL6MaHlgQ98p5bC2bXfSCg2qMI9OMxrrh+W9
rA8HEMLFzqFAbZy2mrflNw37H+u38Y0pSmxJ/fVKTGCzZvRiHJofDHLuZrGL8XvW
KDqFO1VDhel5qIL0333bXaQeft/cDK3OIGFJrjk9S/W6jzdOIevVeQbDoNAc/DqW
jSoM5G4A6dLwYoIEAKqMT9gewl7v88bvSUgZv5gE6A/8yQRqU46eQ7MA12/RM9qy
dK2SjOuANpjjGQpH8PBXJh3+eAGMIHNc+kG54uOVGXwyVgeTfDCIXiFXjK8oRHAF
ROnr21jeA+kFMNEfM/+eHF8JWRiK2lc/6No2cNvgl9rFK1Iavzci6gU7JAwzU6uG
e38SfuwLikn9wnMiD2j6/NSCns1T/pT1YnxGw4qvOW2sTk+xy7dfgXdZbRg4WSSk
`pragma protect end_protected
