	component MebX_Qsys_Project is
		port (
			button_export                                                                                           : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			clk50_clk                                                                                               : in    std_logic                     := 'X';             -- clk
			csense_adc_fo_export                                                                                    : out   std_logic;                                        -- export
			csense_cs_n_export                                                                                      : out   std_logic_vector(1 downto 0);                     -- export
			csense_sck_export                                                                                       : out   std_logic;                                        -- export
			csense_sdi_export                                                                                       : out   std_logic;                                        -- export
			csense_sdo_export                                                                                       : in    std_logic                     := 'X';             -- export
			ctrl_io_lvds_export                                                                                     : out   std_logic_vector(3 downto 0);                     -- export
			dcom_1_sync_end_sync_channel_signal                                                                     : in    std_logic                     := 'X';             -- sync_channel_signal
			dcom_2_sync_end_sync_channel_signal                                                                     : in    std_logic                     := 'X';             -- sync_channel_signal
			dcom_3_sync_end_sync_channel_signal                                                                     : in    std_logic                     := 'X';             -- sync_channel_signal
			dcom_4_sync_end_sync_channel_signal                                                                     : in    std_logic                     := 'X';             -- sync_channel_signal
			dcom_5_sync_end_sync_channel_signal                                                                     : in    std_logic                     := 'X';             -- sync_channel_signal
			dcom_6_sync_end_sync_channel_signal                                                                     : in    std_logic                     := 'X';             -- sync_channel_signal
			dcom_7_sync_end_sync_channel_signal                                                                     : in    std_logic                     := 'X';             -- sync_channel_signal
			dcom_8_sync_end_sync_channel_signal                                                                     : in    std_logic                     := 'X';             -- sync_channel_signal
			dip_export                                                                                              : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			dumb_communication_module_v2_8_conduit_end_rmap_echo_out_echo_en_signal                                 : out   std_logic;                                        -- echo_en_signal
			dumb_communication_module_v2_8_conduit_end_rmap_echo_out_echo_id_en_signal                              : out   std_logic;                                        -- echo_id_en_signal
			dumb_communication_module_v2_8_conduit_end_rmap_echo_out_in_fifo_wrflag_signal                          : out   std_logic;                                        -- in_fifo_wrflag_signal
			dumb_communication_module_v2_8_conduit_end_rmap_echo_out_in_fifo_wrdata_signal                          : out   std_logic_vector(7 downto 0);                     -- in_fifo_wrdata_signal
			dumb_communication_module_v2_8_conduit_end_rmap_echo_out_in_fifo_wrreq_signal                           : out   std_logic;                                        -- in_fifo_wrreq_signal
			dumb_communication_module_v2_8_conduit_end_rmap_echo_out_out_fifo_wrflag_signal                         : out   std_logic;                                        -- out_fifo_wrflag_signal
			dumb_communication_module_v2_8_conduit_end_rmap_echo_out_out_fifo_wrdata_signal                         : out   std_logic_vector(7 downto 0);                     -- out_fifo_wrdata_signal
			dumb_communication_module_v2_8_conduit_end_rmap_echo_out_out_fifo_wrreq_signal                          : out   std_logic;                                        -- out_fifo_wrreq_signal
			dumb_communication_module_v2_timer_avalon_master_data_readdata                                          : in    std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			dumb_communication_module_v2_timer_avalon_master_data_waitrequest                                       : in    std_logic                     := 'X';             -- waitrequest
			dumb_communication_module_v2_timer_avalon_master_data_address                                           : out   std_logic_vector(63 downto 0);                    -- address
			dumb_communication_module_v2_timer_avalon_master_data_read                                              : out   std_logic;                                        -- read
			dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_echo_en_signal                             : out   std_logic;                                        -- echo_en_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_echo_id_en_signal                          : out   std_logic;                                        -- echo_id_en_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_in_fifo_wrflag_signal                      : out   std_logic;                                        -- in_fifo_wrflag_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_in_fifo_wrdata_signal                      : out   std_logic_vector(7 downto 0);                     -- in_fifo_wrdata_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_in_fifo_wrreq_signal                       : out   std_logic;                                        -- in_fifo_wrreq_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_out_fifo_wrflag_signal                     : out   std_logic;                                        -- out_fifo_wrflag_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_out_fifo_wrdata_signal                     : out   std_logic_vector(7 downto 0);                     -- out_fifo_wrdata_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_out_fifo_wrreq_signal                      : out   std_logic;                                        -- out_fifo_wrreq_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_wr_waitrequest_signal                  : in    std_logic                     := 'X';             -- wr_waitrequest_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_readdata_signal                        : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_rd_waitrequest_signal                  : in    std_logic                     := 'X';             -- rd_waitrequest_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_wr_address_signal                      : out   std_logic_vector(31 downto 0);                    -- wr_address_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_write_signal                           : out   std_logic;                                        -- write_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_writedata_signal                       : out   std_logic_vector(7 downto 0);                     -- writedata_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_rd_address_signal                      : out   std_logic_vector(31 downto 0);                    -- rd_address_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_read_signal                            : out   std_logic;                                        -- read_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_mem_configs_out_mem_addr_offset_signal              : out   std_logic_vector(31 downto 0);                    -- mem_addr_offset_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_status_started_signal      : in    std_logic                     := 'X';             -- spw_link_status_started_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_status_connecting_signal   : in    std_logic                     := 'X';             -- spw_link_status_connecting_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_status_running_signal      : in    std_logic                     := 'X';             -- spw_link_status_running_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_error_errdisc_signal       : in    std_logic                     := 'X';             -- spw_link_error_errdisc_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_error_errpar_signal        : in    std_logic                     := 'X';             -- spw_link_error_errpar_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_error_erresc_signal        : in    std_logic                     := 'X';             -- spw_link_error_erresc_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_error_errcred_signal       : in    std_logic                     := 'X';             -- spw_link_error_errcred_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_rx_tick_out_signal     : in    std_logic                     := 'X';             -- spw_timecode_rx_tick_out_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_rx_ctrl_out_signal     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- spw_timecode_rx_ctrl_out_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_rx_time_out_signal     : in    std_logic_vector(5 downto 0)  := (others => 'X'); -- spw_timecode_rx_time_out_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_rx_status_rxvalid_signal   : in    std_logic                     := 'X';             -- spw_data_rx_status_rxvalid_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_rx_status_rxhalff_signal   : in    std_logic                     := 'X';             -- spw_data_rx_status_rxhalff_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_rx_status_rxflag_signal    : in    std_logic                     := 'X';             -- spw_data_rx_status_rxflag_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_rx_status_rxdata_signal    : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- spw_data_rx_status_rxdata_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_tx_status_txrdy_signal     : in    std_logic                     := 'X';             -- spw_data_tx_status_txrdy_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_tx_status_txhalff_signal   : in    std_logic                     := 'X';             -- spw_data_tx_status_txhalff_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_busy_signal  : in    std_logic                     := 'X';             -- spw_errinj_ctrl_errinj_busy_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_ready_signal : in    std_logic                     := 'X';             -- spw_errinj_ctrl_errinj_ready_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_command_enable_signal      : out   std_logic;                                        -- spw_link_command_enable_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_command_autostart_signal   : out   std_logic;                                        -- spw_link_command_autostart_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_command_linkstart_signal   : out   std_logic;                                        -- spw_link_command_linkstart_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_command_linkdis_signal     : out   std_logic;                                        -- spw_link_command_linkdis_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal    : out   std_logic_vector(7 downto 0);                     -- spw_link_command_txdivcnt_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal      : out   std_logic;                                        -- spw_timecode_tx_tick_in_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal      : out   std_logic_vector(1 downto 0);                     -- spw_timecode_tx_ctrl_in_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal      : out   std_logic_vector(5 downto 0);                     -- spw_timecode_tx_time_in_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal   : out   std_logic;                                        -- spw_data_rx_command_rxread_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal  : out   std_logic;                                        -- spw_data_tx_command_txwrite_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal   : out   std_logic;                                        -- spw_data_tx_command_txflag_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal   : out   std_logic_vector(7 downto 0);                     -- spw_data_tx_command_txdata_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_errinj_ctrl_start_errinj_signal : out   std_logic;                                        -- spw_errinj_ctrl_start_errinj_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_errinj_ctrl_reset_errinj_signal : out   std_logic;                                        -- spw_errinj_ctrl_reset_errinj_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_code_signal  : out   std_logic_vector(3 downto 0);                     -- spw_errinj_ctrl_errinj_code_signal
			dumb_communication_module_v2_timer_rprt_interrupt_sender_irq                                            : out   std_logic;                                        -- irq
			dumb_communication_module_v2_timer_sync_conduit_end_sync_channel_signal                                 : in    std_logic                     := 'X';             -- sync_channel_signal
			dumb_communication_module_v2_timer_tx_interrupt_sender_irq                                              : out   std_logic;                                        -- irq
			eth_rst_export                                                                                          : out   std_logic;                                        -- export
			ext_export                                                                                              : in    std_logic                     := 'X';             -- export
			ftdi_clk_clk                                                                                            : in    std_logic                     := 'X';             -- clk
			led_de4_export                                                                                          : out   std_logic_vector(7 downto 0);                     -- export
			led_painel_export                                                                                       : out   std_logic_vector(20 downto 0);                    -- export
			m1_ddr2_i2c_scl_export                                                                                  : out   std_logic;                                        -- export
			m1_ddr2_i2c_sda_export                                                                                  : inout std_logic                     := 'X';             -- export
			m1_ddr2_memory_mem_a                                                                                    : out   std_logic_vector(13 downto 0);                    -- mem_a
			m1_ddr2_memory_mem_ba                                                                                   : out   std_logic_vector(2 downto 0);                     -- mem_ba
			m1_ddr2_memory_mem_ck                                                                                   : out   std_logic_vector(1 downto 0);                     -- mem_ck
			m1_ddr2_memory_mem_ck_n                                                                                 : out   std_logic_vector(1 downto 0);                     -- mem_ck_n
			m1_ddr2_memory_mem_cke                                                                                  : out   std_logic_vector(1 downto 0);                     -- mem_cke
			m1_ddr2_memory_mem_cs_n                                                                                 : out   std_logic_vector(1 downto 0);                     -- mem_cs_n
			m1_ddr2_memory_mem_dm                                                                                   : out   std_logic_vector(7 downto 0);                     -- mem_dm
			m1_ddr2_memory_mem_ras_n                                                                                : out   std_logic_vector(0 downto 0);                     -- mem_ras_n
			m1_ddr2_memory_mem_cas_n                                                                                : out   std_logic_vector(0 downto 0);                     -- mem_cas_n
			m1_ddr2_memory_mem_we_n                                                                                 : out   std_logic_vector(0 downto 0);                     -- mem_we_n
			m1_ddr2_memory_mem_dq                                                                                   : inout std_logic_vector(63 downto 0) := (others => 'X'); -- mem_dq
			m1_ddr2_memory_mem_dqs                                                                                  : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- mem_dqs
			m1_ddr2_memory_mem_dqs_n                                                                                : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- mem_dqs_n
			m1_ddr2_memory_mem_odt                                                                                  : out   std_logic_vector(1 downto 0);                     -- mem_odt
			m1_ddr2_memory_pll_ref_clk_clk                                                                          : in    std_logic                     := 'X';             -- clk
			m1_ddr2_memory_status_local_init_done                                                                   : out   std_logic;                                        -- local_init_done
			m1_ddr2_memory_status_local_cal_success                                                                 : out   std_logic;                                        -- local_cal_success
			m1_ddr2_memory_status_local_cal_fail                                                                    : out   std_logic;                                        -- local_cal_fail
			m1_ddr2_oct_rdn                                                                                         : in    std_logic                     := 'X';             -- rdn
			m1_ddr2_oct_rup                                                                                         : in    std_logic                     := 'X';             -- rup
			m2_ddr2_i2c_scl_export                                                                                  : out   std_logic;                                        -- export
			m2_ddr2_i2c_sda_export                                                                                  : inout std_logic                     := 'X';             -- export
			m2_ddr2_memory_mem_a                                                                                    : out   std_logic_vector(13 downto 0);                    -- mem_a
			m2_ddr2_memory_mem_ba                                                                                   : out   std_logic_vector(2 downto 0);                     -- mem_ba
			m2_ddr2_memory_mem_ck                                                                                   : out   std_logic_vector(1 downto 0);                     -- mem_ck
			m2_ddr2_memory_mem_ck_n                                                                                 : out   std_logic_vector(1 downto 0);                     -- mem_ck_n
			m2_ddr2_memory_mem_cke                                                                                  : out   std_logic_vector(1 downto 0);                     -- mem_cke
			m2_ddr2_memory_mem_cs_n                                                                                 : out   std_logic_vector(1 downto 0);                     -- mem_cs_n
			m2_ddr2_memory_mem_dm                                                                                   : out   std_logic_vector(7 downto 0);                     -- mem_dm
			m2_ddr2_memory_mem_ras_n                                                                                : out   std_logic_vector(0 downto 0);                     -- mem_ras_n
			m2_ddr2_memory_mem_cas_n                                                                                : out   std_logic_vector(0 downto 0);                     -- mem_cas_n
			m2_ddr2_memory_mem_we_n                                                                                 : out   std_logic_vector(0 downto 0);                     -- mem_we_n
			m2_ddr2_memory_mem_dq                                                                                   : inout std_logic_vector(63 downto 0) := (others => 'X'); -- mem_dq
			m2_ddr2_memory_mem_dqs                                                                                  : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- mem_dqs
			m2_ddr2_memory_mem_dqs_n                                                                                : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- mem_dqs_n
			m2_ddr2_memory_mem_odt                                                                                  : out   std_logic_vector(1 downto 0);                     -- mem_odt
			m2_ddr2_memory_dll_sharing_dll_pll_locked                                                               : in    std_logic                     := 'X';             -- dll_pll_locked
			m2_ddr2_memory_dll_sharing_dll_delayctrl                                                                : out   std_logic_vector(5 downto 0);                     -- dll_delayctrl
			m2_ddr2_memory_pll_sharing_pll_mem_clk                                                                  : out   std_logic;                                        -- pll_mem_clk
			m2_ddr2_memory_pll_sharing_pll_write_clk                                                                : out   std_logic;                                        -- pll_write_clk
			m2_ddr2_memory_pll_sharing_pll_locked                                                                   : out   std_logic;                                        -- pll_locked
			m2_ddr2_memory_pll_sharing_pll_write_clk_pre_phy_clk                                                    : out   std_logic;                                        -- pll_write_clk_pre_phy_clk
			m2_ddr2_memory_pll_sharing_pll_addr_cmd_clk                                                             : out   std_logic;                                        -- pll_addr_cmd_clk
			m2_ddr2_memory_pll_sharing_pll_avl_clk                                                                  : out   std_logic;                                        -- pll_avl_clk
			m2_ddr2_memory_pll_sharing_pll_config_clk                                                               : out   std_logic;                                        -- pll_config_clk
			m2_ddr2_memory_status_local_init_done                                                                   : out   std_logic;                                        -- local_init_done
			m2_ddr2_memory_status_local_cal_success                                                                 : out   std_logic;                                        -- local_cal_success
			m2_ddr2_memory_status_local_cal_fail                                                                    : out   std_logic;                                        -- local_cal_fail
			m2_ddr2_oct_rdn                                                                                         : in    std_logic                     := 'X';             -- rdn
			m2_ddr2_oct_rup                                                                                         : in    std_logic                     := 'X';             -- rup
			pio_spw_mux_ch_h_select_export                                                                          : out   std_logic_vector(1 downto 0);                     -- export
			rs232_uart_rxd                                                                                          : in    std_logic                     := 'X';             -- rxd
			rs232_uart_txd                                                                                          : out   std_logic;                                        -- txd
			rst_reset_n                                                                                             : in    std_logic                     := 'X';             -- reset_n
			rst_controller_conduit_reset_input_t_reset_input_signal                                                 : in    std_logic                     := 'X';             -- t_reset_input_signal
			rst_controller_conduit_simucam_reset_t_simucam_reset_signal                                             : out   std_logic;                                        -- t_simucam_reset_signal
			rtcc_alarm_export                                                                                       : in    std_logic                     := 'X';             -- export
			rtcc_cs_n_export                                                                                        : out   std_logic;                                        -- export
			rtcc_sck_export                                                                                         : out   std_logic;                                        -- export
			rtcc_sdi_export                                                                                         : out   std_logic;                                        -- export
			rtcc_sdo_export                                                                                         : in    std_logic                     := 'X';             -- export
			sd_card_ip_b_SD_cmd                                                                                     : inout std_logic                     := 'X';             -- b_SD_cmd
			sd_card_ip_b_SD_dat                                                                                     : inout std_logic                     := 'X';             -- b_SD_dat
			sd_card_ip_b_SD_dat3                                                                                    : inout std_logic                     := 'X';             -- b_SD_dat3
			sd_card_ip_o_SD_clock                                                                                   : out   std_logic;                                        -- o_SD_clock
			sd_card_wp_n_io_export                                                                                  : in    std_logic                     := 'X';             -- export
			spwc_a_enable_spw_rx_enable_signal                                                                      : in    std_logic                     := 'X';             -- spw_rx_enable_signal
			spwc_a_enable_spw_tx_enable_signal                                                                      : in    std_logic                     := 'X';             -- spw_tx_enable_signal
			spwc_a_leds_spw_red_status_led_signal                                                                   : out   std_logic;                                        -- spw_red_status_led_signal
			spwc_a_leds_spw_green_status_led_signal                                                                 : out   std_logic;                                        -- spw_green_status_led_signal
			spwc_a_lvds_spw_lvds_p_data_in_signal                                                                   : in    std_logic                     := 'X';             -- spw_lvds_p_data_in_signal
			spwc_a_lvds_spw_lvds_n_data_in_signal                                                                   : in    std_logic                     := 'X';             -- spw_lvds_n_data_in_signal
			spwc_a_lvds_spw_lvds_p_data_out_signal                                                                  : out   std_logic;                                        -- spw_lvds_p_data_out_signal
			spwc_a_lvds_spw_lvds_n_data_out_signal                                                                  : out   std_logic;                                        -- spw_lvds_n_data_out_signal
			spwc_a_lvds_spw_lvds_p_strobe_out_signal                                                                : out   std_logic;                                        -- spw_lvds_p_strobe_out_signal
			spwc_a_lvds_spw_lvds_n_strobe_out_signal                                                                : out   std_logic;                                        -- spw_lvds_n_strobe_out_signal
			spwc_a_lvds_spw_lvds_p_strobe_in_signal                                                                 : in    std_logic                     := 'X';             -- spw_lvds_p_strobe_in_signal
			spwc_a_lvds_spw_lvds_n_strobe_in_signal                                                                 : in    std_logic                     := 'X';             -- spw_lvds_n_strobe_in_signal
			spwc_b_enable_spw_rx_enable_signal                                                                      : in    std_logic                     := 'X';             -- spw_rx_enable_signal
			spwc_b_enable_spw_tx_enable_signal                                                                      : in    std_logic                     := 'X';             -- spw_tx_enable_signal
			spwc_b_leds_spw_red_status_led_signal                                                                   : out   std_logic;                                        -- spw_red_status_led_signal
			spwc_b_leds_spw_green_status_led_signal                                                                 : out   std_logic;                                        -- spw_green_status_led_signal
			spwc_b_lvds_spw_lvds_p_data_in_signal                                                                   : in    std_logic                     := 'X';             -- spw_lvds_p_data_in_signal
			spwc_b_lvds_spw_lvds_n_data_in_signal                                                                   : in    std_logic                     := 'X';             -- spw_lvds_n_data_in_signal
			spwc_b_lvds_spw_lvds_p_data_out_signal                                                                  : out   std_logic;                                        -- spw_lvds_p_data_out_signal
			spwc_b_lvds_spw_lvds_n_data_out_signal                                                                  : out   std_logic;                                        -- spw_lvds_n_data_out_signal
			spwc_b_lvds_spw_lvds_p_strobe_out_signal                                                                : out   std_logic;                                        -- spw_lvds_p_strobe_out_signal
			spwc_b_lvds_spw_lvds_n_strobe_out_signal                                                                : out   std_logic;                                        -- spw_lvds_n_strobe_out_signal
			spwc_b_lvds_spw_lvds_p_strobe_in_signal                                                                 : in    std_logic                     := 'X';             -- spw_lvds_p_strobe_in_signal
			spwc_b_lvds_spw_lvds_n_strobe_in_signal                                                                 : in    std_logic                     := 'X';             -- spw_lvds_n_strobe_in_signal
			spwc_c_enable_spw_rx_enable_signal                                                                      : in    std_logic                     := 'X';             -- spw_rx_enable_signal
			spwc_c_enable_spw_tx_enable_signal                                                                      : in    std_logic                     := 'X';             -- spw_tx_enable_signal
			spwc_c_leds_spw_red_status_led_signal                                                                   : out   std_logic;                                        -- spw_red_status_led_signal
			spwc_c_leds_spw_green_status_led_signal                                                                 : out   std_logic;                                        -- spw_green_status_led_signal
			spwc_c_lvds_spw_lvds_p_data_in_signal                                                                   : in    std_logic                     := 'X';             -- spw_lvds_p_data_in_signal
			spwc_c_lvds_spw_lvds_n_data_in_signal                                                                   : in    std_logic                     := 'X';             -- spw_lvds_n_data_in_signal
			spwc_c_lvds_spw_lvds_p_data_out_signal                                                                  : out   std_logic;                                        -- spw_lvds_p_data_out_signal
			spwc_c_lvds_spw_lvds_n_data_out_signal                                                                  : out   std_logic;                                        -- spw_lvds_n_data_out_signal
			spwc_c_lvds_spw_lvds_p_strobe_out_signal                                                                : out   std_logic;                                        -- spw_lvds_p_strobe_out_signal
			spwc_c_lvds_spw_lvds_n_strobe_out_signal                                                                : out   std_logic;                                        -- spw_lvds_n_strobe_out_signal
			spwc_c_lvds_spw_lvds_p_strobe_in_signal                                                                 : in    std_logic                     := 'X';             -- spw_lvds_p_strobe_in_signal
			spwc_c_lvds_spw_lvds_n_strobe_in_signal                                                                 : in    std_logic                     := 'X';             -- spw_lvds_n_strobe_in_signal
			spwc_d_enable_spw_rx_enable_signal                                                                      : in    std_logic                     := 'X';             -- spw_rx_enable_signal
			spwc_d_enable_spw_tx_enable_signal                                                                      : in    std_logic                     := 'X';             -- spw_tx_enable_signal
			spwc_d_leds_spw_red_status_led_signal                                                                   : out   std_logic;                                        -- spw_red_status_led_signal
			spwc_d_leds_spw_green_status_led_signal                                                                 : out   std_logic;                                        -- spw_green_status_led_signal
			spwc_d_lvds_spw_lvds_p_data_in_signal                                                                   : in    std_logic                     := 'X';             -- spw_lvds_p_data_in_signal
			spwc_d_lvds_spw_lvds_n_data_in_signal                                                                   : in    std_logic                     := 'X';             -- spw_lvds_n_data_in_signal
			spwc_d_lvds_spw_lvds_p_data_out_signal                                                                  : out   std_logic;                                        -- spw_lvds_p_data_out_signal
			spwc_d_lvds_spw_lvds_n_data_out_signal                                                                  : out   std_logic;                                        -- spw_lvds_n_data_out_signal
			spwc_d_lvds_spw_lvds_p_strobe_out_signal                                                                : out   std_logic;                                        -- spw_lvds_p_strobe_out_signal
			spwc_d_lvds_spw_lvds_n_strobe_out_signal                                                                : out   std_logic;                                        -- spw_lvds_n_strobe_out_signal
			spwc_d_lvds_spw_lvds_p_strobe_in_signal                                                                 : in    std_logic                     := 'X';             -- spw_lvds_p_strobe_in_signal
			spwc_d_lvds_spw_lvds_n_strobe_in_signal                                                                 : in    std_logic                     := 'X';             -- spw_lvds_n_strobe_in_signal
			spwc_e_enable_spw_rx_enable_signal                                                                      : in    std_logic                     := 'X';             -- spw_rx_enable_signal
			spwc_e_enable_spw_tx_enable_signal                                                                      : in    std_logic                     := 'X';             -- spw_tx_enable_signal
			spwc_e_leds_spw_red_status_led_signal                                                                   : out   std_logic;                                        -- spw_red_status_led_signal
			spwc_e_leds_spw_green_status_led_signal                                                                 : out   std_logic;                                        -- spw_green_status_led_signal
			spwc_e_lvds_spw_lvds_p_data_in_signal                                                                   : in    std_logic                     := 'X';             -- spw_lvds_p_data_in_signal
			spwc_e_lvds_spw_lvds_n_data_in_signal                                                                   : in    std_logic                     := 'X';             -- spw_lvds_n_data_in_signal
			spwc_e_lvds_spw_lvds_p_data_out_signal                                                                  : out   std_logic;                                        -- spw_lvds_p_data_out_signal
			spwc_e_lvds_spw_lvds_n_data_out_signal                                                                  : out   std_logic;                                        -- spw_lvds_n_data_out_signal
			spwc_e_lvds_spw_lvds_p_strobe_out_signal                                                                : out   std_logic;                                        -- spw_lvds_p_strobe_out_signal
			spwc_e_lvds_spw_lvds_n_strobe_out_signal                                                                : out   std_logic;                                        -- spw_lvds_n_strobe_out_signal
			spwc_e_lvds_spw_lvds_p_strobe_in_signal                                                                 : in    std_logic                     := 'X';             -- spw_lvds_p_strobe_in_signal
			spwc_e_lvds_spw_lvds_n_strobe_in_signal                                                                 : in    std_logic                     := 'X';             -- spw_lvds_n_strobe_in_signal
			spwc_f_enable_spw_rx_enable_signal                                                                      : in    std_logic                     := 'X';             -- spw_rx_enable_signal
			spwc_f_enable_spw_tx_enable_signal                                                                      : in    std_logic                     := 'X';             -- spw_tx_enable_signal
			spwc_f_leds_spw_red_status_led_signal                                                                   : out   std_logic;                                        -- spw_red_status_led_signal
			spwc_f_leds_spw_green_status_led_signal                                                                 : out   std_logic;                                        -- spw_green_status_led_signal
			spwc_f_lvds_spw_lvds_p_data_in_signal                                                                   : in    std_logic                     := 'X';             -- spw_lvds_p_data_in_signal
			spwc_f_lvds_spw_lvds_n_data_in_signal                                                                   : in    std_logic                     := 'X';             -- spw_lvds_n_data_in_signal
			spwc_f_lvds_spw_lvds_p_data_out_signal                                                                  : out   std_logic;                                        -- spw_lvds_p_data_out_signal
			spwc_f_lvds_spw_lvds_n_data_out_signal                                                                  : out   std_logic;                                        -- spw_lvds_n_data_out_signal
			spwc_f_lvds_spw_lvds_p_strobe_out_signal                                                                : out   std_logic;                                        -- spw_lvds_p_strobe_out_signal
			spwc_f_lvds_spw_lvds_n_strobe_out_signal                                                                : out   std_logic;                                        -- spw_lvds_n_strobe_out_signal
			spwc_f_lvds_spw_lvds_p_strobe_in_signal                                                                 : in    std_logic                     := 'X';             -- spw_lvds_p_strobe_in_signal
			spwc_f_lvds_spw_lvds_n_strobe_in_signal                                                                 : in    std_logic                     := 'X';             -- spw_lvds_n_strobe_in_signal
			spwc_g_enable_spw_rx_enable_signal                                                                      : in    std_logic                     := 'X';             -- spw_rx_enable_signal
			spwc_g_enable_spw_tx_enable_signal                                                                      : in    std_logic                     := 'X';             -- spw_tx_enable_signal
			spwc_g_leds_spw_red_status_led_signal                                                                   : out   std_logic;                                        -- spw_red_status_led_signal
			spwc_g_leds_spw_green_status_led_signal                                                                 : out   std_logic;                                        -- spw_green_status_led_signal
			spwc_g_lvds_spw_lvds_p_data_in_signal                                                                   : in    std_logic                     := 'X';             -- spw_lvds_p_data_in_signal
			spwc_g_lvds_spw_lvds_n_data_in_signal                                                                   : in    std_logic                     := 'X';             -- spw_lvds_n_data_in_signal
			spwc_g_lvds_spw_lvds_p_data_out_signal                                                                  : out   std_logic;                                        -- spw_lvds_p_data_out_signal
			spwc_g_lvds_spw_lvds_n_data_out_signal                                                                  : out   std_logic;                                        -- spw_lvds_n_data_out_signal
			spwc_g_lvds_spw_lvds_p_strobe_out_signal                                                                : out   std_logic;                                        -- spw_lvds_p_strobe_out_signal
			spwc_g_lvds_spw_lvds_n_strobe_out_signal                                                                : out   std_logic;                                        -- spw_lvds_n_strobe_out_signal
			spwc_g_lvds_spw_lvds_p_strobe_in_signal                                                                 : in    std_logic                     := 'X';             -- spw_lvds_p_strobe_in_signal
			spwc_g_lvds_spw_lvds_n_strobe_in_signal                                                                 : in    std_logic                     := 'X';             -- spw_lvds_n_strobe_in_signal
			spwc_h_enable_spw_rx_enable_signal                                                                      : in    std_logic                     := 'X';             -- spw_rx_enable_signal
			spwc_h_enable_spw_tx_enable_signal                                                                      : in    std_logic                     := 'X';             -- spw_tx_enable_signal
			spwc_h_leds_spw_red_status_led_signal                                                                   : out   std_logic;                                        -- spw_red_status_led_signal
			spwc_h_leds_spw_green_status_led_signal                                                                 : out   std_logic;                                        -- spw_green_status_led_signal
			spwc_h_lvds_spw_lvds_p_data_in_signal                                                                   : in    std_logic                     := 'X';             -- spw_lvds_p_data_in_signal
			spwc_h_lvds_spw_lvds_n_data_in_signal                                                                   : in    std_logic                     := 'X';             -- spw_lvds_n_data_in_signal
			spwc_h_lvds_spw_lvds_p_data_out_signal                                                                  : out   std_logic;                                        -- spw_lvds_p_data_out_signal
			spwc_h_lvds_spw_lvds_n_data_out_signal                                                                  : out   std_logic;                                        -- spw_lvds_n_data_out_signal
			spwc_h_lvds_spw_lvds_p_strobe_out_signal                                                                : out   std_logic;                                        -- spw_lvds_p_strobe_out_signal
			spwc_h_lvds_spw_lvds_n_strobe_out_signal                                                                : out   std_logic;                                        -- spw_lvds_n_strobe_out_signal
			spwc_h_lvds_spw_lvds_p_strobe_in_signal                                                                 : in    std_logic                     := 'X';             -- spw_lvds_p_strobe_in_signal
			spwc_h_lvds_spw_lvds_n_strobe_in_signal                                                                 : in    std_logic                     := 'X';             -- spw_lvds_n_strobe_in_signal
			spwm_h_select_mux_select_signal                                                                         : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- mux_select_signal
			ssdp_ssdp0                                                                                              : out   std_logic_vector(7 downto 0);                     -- ssdp0
			ssdp_ssdp1                                                                                              : out   std_logic_vector(7 downto 0);                     -- ssdp1
			sync_in_conduit                                                                                         : in    std_logic                     := 'X';             -- conduit
			sync_in_en_conduit                                                                                      : in    std_logic                     := 'X';             -- conduit
			sync_out_conduit                                                                                        : out   std_logic;                                        -- conduit
			sync_out_en_conduit                                                                                     : in    std_logic                     := 'X';             -- conduit
			sync_spw1_conduit                                                                                       : out   std_logic;                                        -- conduit
			sync_spw2_conduit                                                                                       : out   std_logic;                                        -- conduit
			sync_spw3_conduit                                                                                       : out   std_logic;                                        -- conduit
			sync_spw4_conduit                                                                                       : out   std_logic;                                        -- conduit
			sync_spw5_conduit                                                                                       : out   std_logic;                                        -- conduit
			sync_spw6_conduit                                                                                       : out   std_logic;                                        -- conduit
			sync_spw7_conduit                                                                                       : out   std_logic;                                        -- conduit
			sync_spw8_conduit                                                                                       : out   std_logic;                                        -- conduit
			temp_scl_export                                                                                         : out   std_logic;                                        -- export
			temp_sda_export                                                                                         : inout std_logic                     := 'X';             -- export
			timer_1ms_external_port_export                                                                          : out   std_logic;                                        -- export
			timer_1us_external_port_export                                                                          : out   std_logic;                                        -- export
			tristate_conduit_tcm_address_out                                                                        : out   std_logic_vector(25 downto 0);                    -- tcm_address_out
			tristate_conduit_tcm_read_n_out                                                                         : out   std_logic_vector(0 downto 0);                     -- tcm_read_n_out
			tristate_conduit_tcm_write_n_out                                                                        : out   std_logic_vector(0 downto 0);                     -- tcm_write_n_out
			tristate_conduit_tcm_data_out                                                                           : inout std_logic_vector(15 downto 0) := (others => 'X'); -- tcm_data_out
			tristate_conduit_tcm_chipselect_n_out                                                                   : out   std_logic_vector(0 downto 0);                     -- tcm_chipselect_n_out
			umft601a_pins_umft_clock_signal                                                                         : in    std_logic                     := 'X';             -- umft_clock_signal
			umft601a_pins_umft_txe_n_signal                                                                         : in    std_logic                     := 'X';             -- umft_txe_n_signal
			umft601a_pins_umft_rxf_n_signal                                                                         : in    std_logic                     := 'X';             -- umft_rxf_n_signal
			umft601a_pins_umft_data_signal                                                                          : inout std_logic_vector(31 downto 0) := (others => 'X'); -- umft_data_signal
			umft601a_pins_umft_be_signal                                                                            : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- umft_be_signal
			umft601a_pins_umft_wakeup_n_signal                                                                      : inout std_logic                     := 'X';             -- umft_wakeup_n_signal
			umft601a_pins_umft_gpio_bus_signal                                                                      : inout std_logic_vector(1 downto 0)  := (others => 'X'); -- umft_gpio_bus_signal
			umft601a_pins_umft_reset_n_signal                                                                       : out   std_logic;                                        -- umft_reset_n_signal
			umft601a_pins_umft_wr_n_signal                                                                          : out   std_logic;                                        -- umft_wr_n_signal
			umft601a_pins_umft_rd_n_signal                                                                          : out   std_logic;                                        -- umft_rd_n_signal
			umft601a_pins_umft_oe_n_signal                                                                          : out   std_logic;                                        -- umft_oe_n_signal
			umft601a_pins_umft_siwu_n_signal                                                                        : out   std_logic                                         -- umft_siwu_n_signal
		);
	end component MebX_Qsys_Project;

	u0 : component MebX_Qsys_Project
		port map (
			button_export                                                                                           => CONNECTED_TO_button_export,                                                                                           --                                                              button.export
			clk50_clk                                                                                               => CONNECTED_TO_clk50_clk,                                                                                               --                                                               clk50.clk
			csense_adc_fo_export                                                                                    => CONNECTED_TO_csense_adc_fo_export,                                                                                    --                                                       csense_adc_fo.export
			csense_cs_n_export                                                                                      => CONNECTED_TO_csense_cs_n_export,                                                                                      --                                                         csense_cs_n.export
			csense_sck_export                                                                                       => CONNECTED_TO_csense_sck_export,                                                                                       --                                                          csense_sck.export
			csense_sdi_export                                                                                       => CONNECTED_TO_csense_sdi_export,                                                                                       --                                                          csense_sdi.export
			csense_sdo_export                                                                                       => CONNECTED_TO_csense_sdo_export,                                                                                       --                                                          csense_sdo.export
			ctrl_io_lvds_export                                                                                     => CONNECTED_TO_ctrl_io_lvds_export,                                                                                     --                                                        ctrl_io_lvds.export
			dcom_1_sync_end_sync_channel_signal                                                                     => CONNECTED_TO_dcom_1_sync_end_sync_channel_signal,                                                                     --                                                     dcom_1_sync_end.sync_channel_signal
			dcom_2_sync_end_sync_channel_signal                                                                     => CONNECTED_TO_dcom_2_sync_end_sync_channel_signal,                                                                     --                                                     dcom_2_sync_end.sync_channel_signal
			dcom_3_sync_end_sync_channel_signal                                                                     => CONNECTED_TO_dcom_3_sync_end_sync_channel_signal,                                                                     --                                                     dcom_3_sync_end.sync_channel_signal
			dcom_4_sync_end_sync_channel_signal                                                                     => CONNECTED_TO_dcom_4_sync_end_sync_channel_signal,                                                                     --                                                     dcom_4_sync_end.sync_channel_signal
			dcom_5_sync_end_sync_channel_signal                                                                     => CONNECTED_TO_dcom_5_sync_end_sync_channel_signal,                                                                     --                                                     dcom_5_sync_end.sync_channel_signal
			dcom_6_sync_end_sync_channel_signal                                                                     => CONNECTED_TO_dcom_6_sync_end_sync_channel_signal,                                                                     --                                                     dcom_6_sync_end.sync_channel_signal
			dcom_7_sync_end_sync_channel_signal                                                                     => CONNECTED_TO_dcom_7_sync_end_sync_channel_signal,                                                                     --                                                     dcom_7_sync_end.sync_channel_signal
			dcom_8_sync_end_sync_channel_signal                                                                     => CONNECTED_TO_dcom_8_sync_end_sync_channel_signal,                                                                     --                                                     dcom_8_sync_end.sync_channel_signal
			dip_export                                                                                              => CONNECTED_TO_dip_export,                                                                                              --                                                                 dip.export
			dumb_communication_module_v2_8_conduit_end_rmap_echo_out_echo_en_signal                                 => CONNECTED_TO_dumb_communication_module_v2_8_conduit_end_rmap_echo_out_echo_en_signal,                                 --            dumb_communication_module_v2_8_conduit_end_rmap_echo_out.echo_en_signal
			dumb_communication_module_v2_8_conduit_end_rmap_echo_out_echo_id_en_signal                              => CONNECTED_TO_dumb_communication_module_v2_8_conduit_end_rmap_echo_out_echo_id_en_signal,                              --                                                                    .echo_id_en_signal
			dumb_communication_module_v2_8_conduit_end_rmap_echo_out_in_fifo_wrflag_signal                          => CONNECTED_TO_dumb_communication_module_v2_8_conduit_end_rmap_echo_out_in_fifo_wrflag_signal,                          --                                                                    .in_fifo_wrflag_signal
			dumb_communication_module_v2_8_conduit_end_rmap_echo_out_in_fifo_wrdata_signal                          => CONNECTED_TO_dumb_communication_module_v2_8_conduit_end_rmap_echo_out_in_fifo_wrdata_signal,                          --                                                                    .in_fifo_wrdata_signal
			dumb_communication_module_v2_8_conduit_end_rmap_echo_out_in_fifo_wrreq_signal                           => CONNECTED_TO_dumb_communication_module_v2_8_conduit_end_rmap_echo_out_in_fifo_wrreq_signal,                           --                                                                    .in_fifo_wrreq_signal
			dumb_communication_module_v2_8_conduit_end_rmap_echo_out_out_fifo_wrflag_signal                         => CONNECTED_TO_dumb_communication_module_v2_8_conduit_end_rmap_echo_out_out_fifo_wrflag_signal,                         --                                                                    .out_fifo_wrflag_signal
			dumb_communication_module_v2_8_conduit_end_rmap_echo_out_out_fifo_wrdata_signal                         => CONNECTED_TO_dumb_communication_module_v2_8_conduit_end_rmap_echo_out_out_fifo_wrdata_signal,                         --                                                                    .out_fifo_wrdata_signal
			dumb_communication_module_v2_8_conduit_end_rmap_echo_out_out_fifo_wrreq_signal                          => CONNECTED_TO_dumb_communication_module_v2_8_conduit_end_rmap_echo_out_out_fifo_wrreq_signal,                          --                                                                    .out_fifo_wrreq_signal
			dumb_communication_module_v2_timer_avalon_master_data_readdata                                          => CONNECTED_TO_dumb_communication_module_v2_timer_avalon_master_data_readdata,                                          --               dumb_communication_module_v2_timer_avalon_master_data.readdata
			dumb_communication_module_v2_timer_avalon_master_data_waitrequest                                       => CONNECTED_TO_dumb_communication_module_v2_timer_avalon_master_data_waitrequest,                                       --                                                                    .waitrequest
			dumb_communication_module_v2_timer_avalon_master_data_address                                           => CONNECTED_TO_dumb_communication_module_v2_timer_avalon_master_data_address,                                           --                                                                    .address
			dumb_communication_module_v2_timer_avalon_master_data_read                                              => CONNECTED_TO_dumb_communication_module_v2_timer_avalon_master_data_read,                                              --                                                                    .read
			dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_echo_en_signal                             => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_echo_en_signal,                             --        dumb_communication_module_v2_timer_conduit_end_rmap_echo_out.echo_en_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_echo_id_en_signal                          => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_echo_id_en_signal,                          --                                                                    .echo_id_en_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_in_fifo_wrflag_signal                      => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_in_fifo_wrflag_signal,                      --                                                                    .in_fifo_wrflag_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_in_fifo_wrdata_signal                      => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_in_fifo_wrdata_signal,                      --                                                                    .in_fifo_wrdata_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_in_fifo_wrreq_signal                       => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_in_fifo_wrreq_signal,                       --                                                                    .in_fifo_wrreq_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_out_fifo_wrflag_signal                     => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_out_fifo_wrflag_signal,                     --                                                                    .out_fifo_wrflag_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_out_fifo_wrdata_signal                     => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_out_fifo_wrdata_signal,                     --                                                                    .out_fifo_wrdata_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_out_fifo_wrreq_signal                      => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_echo_out_out_fifo_wrreq_signal,                      --                                                                    .out_fifo_wrreq_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_wr_waitrequest_signal                  => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_wr_waitrequest_signal,                  --    dumb_communication_module_v2_timer_conduit_end_rmap_master_codec.wr_waitrequest_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_readdata_signal                        => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_readdata_signal,                        --                                                                    .readdata_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_rd_waitrequest_signal                  => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_rd_waitrequest_signal,                  --                                                                    .rd_waitrequest_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_wr_address_signal                      => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_wr_address_signal,                      --                                                                    .wr_address_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_write_signal                           => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_write_signal,                           --                                                                    .write_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_writedata_signal                       => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_writedata_signal,                       --                                                                    .writedata_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_rd_address_signal                      => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_rd_address_signal,                      --                                                                    .rd_address_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_read_signal                            => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_master_codec_read_signal,                            --                                                                    .read_signal
			dumb_communication_module_v2_timer_conduit_end_rmap_mem_configs_out_mem_addr_offset_signal              => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_rmap_mem_configs_out_mem_addr_offset_signal,              -- dumb_communication_module_v2_timer_conduit_end_rmap_mem_configs_out.mem_addr_offset_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_status_started_signal      => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_status_started_signal,      -- dumb_communication_module_v2_timer_conduit_end_spacewire_controller.spw_link_status_started_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_status_connecting_signal   => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_status_connecting_signal,   --                                                                    .spw_link_status_connecting_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_status_running_signal      => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_status_running_signal,      --                                                                    .spw_link_status_running_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_error_errdisc_signal       => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_error_errdisc_signal,       --                                                                    .spw_link_error_errdisc_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_error_errpar_signal        => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_error_errpar_signal,        --                                                                    .spw_link_error_errpar_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_error_erresc_signal        => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_error_erresc_signal,        --                                                                    .spw_link_error_erresc_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_error_errcred_signal       => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_error_errcred_signal,       --                                                                    .spw_link_error_errcred_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_rx_tick_out_signal     => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_rx_tick_out_signal,     --                                                                    .spw_timecode_rx_tick_out_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_rx_ctrl_out_signal     => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_rx_ctrl_out_signal,     --                                                                    .spw_timecode_rx_ctrl_out_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_rx_time_out_signal     => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_rx_time_out_signal,     --                                                                    .spw_timecode_rx_time_out_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_rx_status_rxvalid_signal   => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_rx_status_rxvalid_signal,   --                                                                    .spw_data_rx_status_rxvalid_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_rx_status_rxhalff_signal   => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_rx_status_rxhalff_signal,   --                                                                    .spw_data_rx_status_rxhalff_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_rx_status_rxflag_signal    => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_rx_status_rxflag_signal,    --                                                                    .spw_data_rx_status_rxflag_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_rx_status_rxdata_signal    => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_rx_status_rxdata_signal,    --                                                                    .spw_data_rx_status_rxdata_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_tx_status_txrdy_signal     => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_tx_status_txrdy_signal,     --                                                                    .spw_data_tx_status_txrdy_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_tx_status_txhalff_signal   => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_tx_status_txhalff_signal,   --                                                                    .spw_data_tx_status_txhalff_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_busy_signal  => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_busy_signal,  --                                                                    .spw_errinj_ctrl_errinj_busy_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_ready_signal => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_ready_signal, --                                                                    .spw_errinj_ctrl_errinj_ready_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_command_enable_signal      => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_command_enable_signal,      --                                                                    .spw_link_command_enable_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_command_autostart_signal   => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_command_autostart_signal,   --                                                                    .spw_link_command_autostart_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_command_linkstart_signal   => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_command_linkstart_signal,   --                                                                    .spw_link_command_linkstart_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_command_linkdis_signal     => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_command_linkdis_signal,     --                                                                    .spw_link_command_linkdis_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal    => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal,    --                                                                    .spw_link_command_txdivcnt_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal      => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal,      --                                                                    .spw_timecode_tx_tick_in_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal      => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal,      --                                                                    .spw_timecode_tx_ctrl_in_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal      => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal,      --                                                                    .spw_timecode_tx_time_in_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal   => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal,   --                                                                    .spw_data_rx_command_rxread_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal  => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal,  --                                                                    .spw_data_tx_command_txwrite_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal   => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal,   --                                                                    .spw_data_tx_command_txflag_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal   => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal,   --                                                                    .spw_data_tx_command_txdata_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_errinj_ctrl_start_errinj_signal => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_errinj_ctrl_start_errinj_signal, --                                                                    .spw_errinj_ctrl_start_errinj_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_errinj_ctrl_reset_errinj_signal => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_errinj_ctrl_reset_errinj_signal, --                                                                    .spw_errinj_ctrl_reset_errinj_signal
			dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_code_signal  => CONNECTED_TO_dumb_communication_module_v2_timer_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_code_signal,  --                                                                    .spw_errinj_ctrl_errinj_code_signal
			dumb_communication_module_v2_timer_rprt_interrupt_sender_irq                                            => CONNECTED_TO_dumb_communication_module_v2_timer_rprt_interrupt_sender_irq,                                            --            dumb_communication_module_v2_timer_rprt_interrupt_sender.irq
			dumb_communication_module_v2_timer_sync_conduit_end_sync_channel_signal                                 => CONNECTED_TO_dumb_communication_module_v2_timer_sync_conduit_end_sync_channel_signal,                                 --                 dumb_communication_module_v2_timer_sync_conduit_end.sync_channel_signal
			dumb_communication_module_v2_timer_tx_interrupt_sender_irq                                              => CONNECTED_TO_dumb_communication_module_v2_timer_tx_interrupt_sender_irq,                                              --              dumb_communication_module_v2_timer_tx_interrupt_sender.irq
			eth_rst_export                                                                                          => CONNECTED_TO_eth_rst_export,                                                                                          --                                                             eth_rst.export
			ext_export                                                                                              => CONNECTED_TO_ext_export,                                                                                              --                                                                 ext.export
			ftdi_clk_clk                                                                                            => CONNECTED_TO_ftdi_clk_clk,                                                                                            --                                                            ftdi_clk.clk
			led_de4_export                                                                                          => CONNECTED_TO_led_de4_export,                                                                                          --                                                             led_de4.export
			led_painel_export                                                                                       => CONNECTED_TO_led_painel_export,                                                                                       --                                                          led_painel.export
			m1_ddr2_i2c_scl_export                                                                                  => CONNECTED_TO_m1_ddr2_i2c_scl_export,                                                                                  --                                                     m1_ddr2_i2c_scl.export
			m1_ddr2_i2c_sda_export                                                                                  => CONNECTED_TO_m1_ddr2_i2c_sda_export,                                                                                  --                                                     m1_ddr2_i2c_sda.export
			m1_ddr2_memory_mem_a                                                                                    => CONNECTED_TO_m1_ddr2_memory_mem_a,                                                                                    --                                                      m1_ddr2_memory.mem_a
			m1_ddr2_memory_mem_ba                                                                                   => CONNECTED_TO_m1_ddr2_memory_mem_ba,                                                                                   --                                                                    .mem_ba
			m1_ddr2_memory_mem_ck                                                                                   => CONNECTED_TO_m1_ddr2_memory_mem_ck,                                                                                   --                                                                    .mem_ck
			m1_ddr2_memory_mem_ck_n                                                                                 => CONNECTED_TO_m1_ddr2_memory_mem_ck_n,                                                                                 --                                                                    .mem_ck_n
			m1_ddr2_memory_mem_cke                                                                                  => CONNECTED_TO_m1_ddr2_memory_mem_cke,                                                                                  --                                                                    .mem_cke
			m1_ddr2_memory_mem_cs_n                                                                                 => CONNECTED_TO_m1_ddr2_memory_mem_cs_n,                                                                                 --                                                                    .mem_cs_n
			m1_ddr2_memory_mem_dm                                                                                   => CONNECTED_TO_m1_ddr2_memory_mem_dm,                                                                                   --                                                                    .mem_dm
			m1_ddr2_memory_mem_ras_n                                                                                => CONNECTED_TO_m1_ddr2_memory_mem_ras_n,                                                                                --                                                                    .mem_ras_n
			m1_ddr2_memory_mem_cas_n                                                                                => CONNECTED_TO_m1_ddr2_memory_mem_cas_n,                                                                                --                                                                    .mem_cas_n
			m1_ddr2_memory_mem_we_n                                                                                 => CONNECTED_TO_m1_ddr2_memory_mem_we_n,                                                                                 --                                                                    .mem_we_n
			m1_ddr2_memory_mem_dq                                                                                   => CONNECTED_TO_m1_ddr2_memory_mem_dq,                                                                                   --                                                                    .mem_dq
			m1_ddr2_memory_mem_dqs                                                                                  => CONNECTED_TO_m1_ddr2_memory_mem_dqs,                                                                                  --                                                                    .mem_dqs
			m1_ddr2_memory_mem_dqs_n                                                                                => CONNECTED_TO_m1_ddr2_memory_mem_dqs_n,                                                                                --                                                                    .mem_dqs_n
			m1_ddr2_memory_mem_odt                                                                                  => CONNECTED_TO_m1_ddr2_memory_mem_odt,                                                                                  --                                                                    .mem_odt
			m1_ddr2_memory_pll_ref_clk_clk                                                                          => CONNECTED_TO_m1_ddr2_memory_pll_ref_clk_clk,                                                                          --                                          m1_ddr2_memory_pll_ref_clk.clk
			m1_ddr2_memory_status_local_init_done                                                                   => CONNECTED_TO_m1_ddr2_memory_status_local_init_done,                                                                   --                                               m1_ddr2_memory_status.local_init_done
			m1_ddr2_memory_status_local_cal_success                                                                 => CONNECTED_TO_m1_ddr2_memory_status_local_cal_success,                                                                 --                                                                    .local_cal_success
			m1_ddr2_memory_status_local_cal_fail                                                                    => CONNECTED_TO_m1_ddr2_memory_status_local_cal_fail,                                                                    --                                                                    .local_cal_fail
			m1_ddr2_oct_rdn                                                                                         => CONNECTED_TO_m1_ddr2_oct_rdn,                                                                                         --                                                         m1_ddr2_oct.rdn
			m1_ddr2_oct_rup                                                                                         => CONNECTED_TO_m1_ddr2_oct_rup,                                                                                         --                                                                    .rup
			m2_ddr2_i2c_scl_export                                                                                  => CONNECTED_TO_m2_ddr2_i2c_scl_export,                                                                                  --                                                     m2_ddr2_i2c_scl.export
			m2_ddr2_i2c_sda_export                                                                                  => CONNECTED_TO_m2_ddr2_i2c_sda_export,                                                                                  --                                                     m2_ddr2_i2c_sda.export
			m2_ddr2_memory_mem_a                                                                                    => CONNECTED_TO_m2_ddr2_memory_mem_a,                                                                                    --                                                      m2_ddr2_memory.mem_a
			m2_ddr2_memory_mem_ba                                                                                   => CONNECTED_TO_m2_ddr2_memory_mem_ba,                                                                                   --                                                                    .mem_ba
			m2_ddr2_memory_mem_ck                                                                                   => CONNECTED_TO_m2_ddr2_memory_mem_ck,                                                                                   --                                                                    .mem_ck
			m2_ddr2_memory_mem_ck_n                                                                                 => CONNECTED_TO_m2_ddr2_memory_mem_ck_n,                                                                                 --                                                                    .mem_ck_n
			m2_ddr2_memory_mem_cke                                                                                  => CONNECTED_TO_m2_ddr2_memory_mem_cke,                                                                                  --                                                                    .mem_cke
			m2_ddr2_memory_mem_cs_n                                                                                 => CONNECTED_TO_m2_ddr2_memory_mem_cs_n,                                                                                 --                                                                    .mem_cs_n
			m2_ddr2_memory_mem_dm                                                                                   => CONNECTED_TO_m2_ddr2_memory_mem_dm,                                                                                   --                                                                    .mem_dm
			m2_ddr2_memory_mem_ras_n                                                                                => CONNECTED_TO_m2_ddr2_memory_mem_ras_n,                                                                                --                                                                    .mem_ras_n
			m2_ddr2_memory_mem_cas_n                                                                                => CONNECTED_TO_m2_ddr2_memory_mem_cas_n,                                                                                --                                                                    .mem_cas_n
			m2_ddr2_memory_mem_we_n                                                                                 => CONNECTED_TO_m2_ddr2_memory_mem_we_n,                                                                                 --                                                                    .mem_we_n
			m2_ddr2_memory_mem_dq                                                                                   => CONNECTED_TO_m2_ddr2_memory_mem_dq,                                                                                   --                                                                    .mem_dq
			m2_ddr2_memory_mem_dqs                                                                                  => CONNECTED_TO_m2_ddr2_memory_mem_dqs,                                                                                  --                                                                    .mem_dqs
			m2_ddr2_memory_mem_dqs_n                                                                                => CONNECTED_TO_m2_ddr2_memory_mem_dqs_n,                                                                                --                                                                    .mem_dqs_n
			m2_ddr2_memory_mem_odt                                                                                  => CONNECTED_TO_m2_ddr2_memory_mem_odt,                                                                                  --                                                                    .mem_odt
			m2_ddr2_memory_dll_sharing_dll_pll_locked                                                               => CONNECTED_TO_m2_ddr2_memory_dll_sharing_dll_pll_locked,                                                               --                                          m2_ddr2_memory_dll_sharing.dll_pll_locked
			m2_ddr2_memory_dll_sharing_dll_delayctrl                                                                => CONNECTED_TO_m2_ddr2_memory_dll_sharing_dll_delayctrl,                                                                --                                                                    .dll_delayctrl
			m2_ddr2_memory_pll_sharing_pll_mem_clk                                                                  => CONNECTED_TO_m2_ddr2_memory_pll_sharing_pll_mem_clk,                                                                  --                                          m2_ddr2_memory_pll_sharing.pll_mem_clk
			m2_ddr2_memory_pll_sharing_pll_write_clk                                                                => CONNECTED_TO_m2_ddr2_memory_pll_sharing_pll_write_clk,                                                                --                                                                    .pll_write_clk
			m2_ddr2_memory_pll_sharing_pll_locked                                                                   => CONNECTED_TO_m2_ddr2_memory_pll_sharing_pll_locked,                                                                   --                                                                    .pll_locked
			m2_ddr2_memory_pll_sharing_pll_write_clk_pre_phy_clk                                                    => CONNECTED_TO_m2_ddr2_memory_pll_sharing_pll_write_clk_pre_phy_clk,                                                    --                                                                    .pll_write_clk_pre_phy_clk
			m2_ddr2_memory_pll_sharing_pll_addr_cmd_clk                                                             => CONNECTED_TO_m2_ddr2_memory_pll_sharing_pll_addr_cmd_clk,                                                             --                                                                    .pll_addr_cmd_clk
			m2_ddr2_memory_pll_sharing_pll_avl_clk                                                                  => CONNECTED_TO_m2_ddr2_memory_pll_sharing_pll_avl_clk,                                                                  --                                                                    .pll_avl_clk
			m2_ddr2_memory_pll_sharing_pll_config_clk                                                               => CONNECTED_TO_m2_ddr2_memory_pll_sharing_pll_config_clk,                                                               --                                                                    .pll_config_clk
			m2_ddr2_memory_status_local_init_done                                                                   => CONNECTED_TO_m2_ddr2_memory_status_local_init_done,                                                                   --                                               m2_ddr2_memory_status.local_init_done
			m2_ddr2_memory_status_local_cal_success                                                                 => CONNECTED_TO_m2_ddr2_memory_status_local_cal_success,                                                                 --                                                                    .local_cal_success
			m2_ddr2_memory_status_local_cal_fail                                                                    => CONNECTED_TO_m2_ddr2_memory_status_local_cal_fail,                                                                    --                                                                    .local_cal_fail
			m2_ddr2_oct_rdn                                                                                         => CONNECTED_TO_m2_ddr2_oct_rdn,                                                                                         --                                                         m2_ddr2_oct.rdn
			m2_ddr2_oct_rup                                                                                         => CONNECTED_TO_m2_ddr2_oct_rup,                                                                                         --                                                                    .rup
			pio_spw_mux_ch_h_select_export                                                                          => CONNECTED_TO_pio_spw_mux_ch_h_select_export,                                                                          --                                             pio_spw_mux_ch_h_select.export
			rs232_uart_rxd                                                                                          => CONNECTED_TO_rs232_uart_rxd,                                                                                          --                                                          rs232_uart.rxd
			rs232_uart_txd                                                                                          => CONNECTED_TO_rs232_uart_txd,                                                                                          --                                                                    .txd
			rst_reset_n                                                                                             => CONNECTED_TO_rst_reset_n,                                                                                             --                                                                 rst.reset_n
			rst_controller_conduit_reset_input_t_reset_input_signal                                                 => CONNECTED_TO_rst_controller_conduit_reset_input_t_reset_input_signal,                                                 --                                  rst_controller_conduit_reset_input.t_reset_input_signal
			rst_controller_conduit_simucam_reset_t_simucam_reset_signal                                             => CONNECTED_TO_rst_controller_conduit_simucam_reset_t_simucam_reset_signal,                                             --                                rst_controller_conduit_simucam_reset.t_simucam_reset_signal
			rtcc_alarm_export                                                                                       => CONNECTED_TO_rtcc_alarm_export,                                                                                       --                                                          rtcc_alarm.export
			rtcc_cs_n_export                                                                                        => CONNECTED_TO_rtcc_cs_n_export,                                                                                        --                                                           rtcc_cs_n.export
			rtcc_sck_export                                                                                         => CONNECTED_TO_rtcc_sck_export,                                                                                         --                                                            rtcc_sck.export
			rtcc_sdi_export                                                                                         => CONNECTED_TO_rtcc_sdi_export,                                                                                         --                                                            rtcc_sdi.export
			rtcc_sdo_export                                                                                         => CONNECTED_TO_rtcc_sdo_export,                                                                                         --                                                            rtcc_sdo.export
			sd_card_ip_b_SD_cmd                                                                                     => CONNECTED_TO_sd_card_ip_b_SD_cmd,                                                                                     --                                                          sd_card_ip.b_SD_cmd
			sd_card_ip_b_SD_dat                                                                                     => CONNECTED_TO_sd_card_ip_b_SD_dat,                                                                                     --                                                                    .b_SD_dat
			sd_card_ip_b_SD_dat3                                                                                    => CONNECTED_TO_sd_card_ip_b_SD_dat3,                                                                                    --                                                                    .b_SD_dat3
			sd_card_ip_o_SD_clock                                                                                   => CONNECTED_TO_sd_card_ip_o_SD_clock,                                                                                   --                                                                    .o_SD_clock
			sd_card_wp_n_io_export                                                                                  => CONNECTED_TO_sd_card_wp_n_io_export,                                                                                  --                                                     sd_card_wp_n_io.export
			spwc_a_enable_spw_rx_enable_signal                                                                      => CONNECTED_TO_spwc_a_enable_spw_rx_enable_signal,                                                                      --                                                       spwc_a_enable.spw_rx_enable_signal
			spwc_a_enable_spw_tx_enable_signal                                                                      => CONNECTED_TO_spwc_a_enable_spw_tx_enable_signal,                                                                      --                                                                    .spw_tx_enable_signal
			spwc_a_leds_spw_red_status_led_signal                                                                   => CONNECTED_TO_spwc_a_leds_spw_red_status_led_signal,                                                                   --                                                         spwc_a_leds.spw_red_status_led_signal
			spwc_a_leds_spw_green_status_led_signal                                                                 => CONNECTED_TO_spwc_a_leds_spw_green_status_led_signal,                                                                 --                                                                    .spw_green_status_led_signal
			spwc_a_lvds_spw_lvds_p_data_in_signal                                                                   => CONNECTED_TO_spwc_a_lvds_spw_lvds_p_data_in_signal,                                                                   --                                                         spwc_a_lvds.spw_lvds_p_data_in_signal
			spwc_a_lvds_spw_lvds_n_data_in_signal                                                                   => CONNECTED_TO_spwc_a_lvds_spw_lvds_n_data_in_signal,                                                                   --                                                                    .spw_lvds_n_data_in_signal
			spwc_a_lvds_spw_lvds_p_data_out_signal                                                                  => CONNECTED_TO_spwc_a_lvds_spw_lvds_p_data_out_signal,                                                                  --                                                                    .spw_lvds_p_data_out_signal
			spwc_a_lvds_spw_lvds_n_data_out_signal                                                                  => CONNECTED_TO_spwc_a_lvds_spw_lvds_n_data_out_signal,                                                                  --                                                                    .spw_lvds_n_data_out_signal
			spwc_a_lvds_spw_lvds_p_strobe_out_signal                                                                => CONNECTED_TO_spwc_a_lvds_spw_lvds_p_strobe_out_signal,                                                                --                                                                    .spw_lvds_p_strobe_out_signal
			spwc_a_lvds_spw_lvds_n_strobe_out_signal                                                                => CONNECTED_TO_spwc_a_lvds_spw_lvds_n_strobe_out_signal,                                                                --                                                                    .spw_lvds_n_strobe_out_signal
			spwc_a_lvds_spw_lvds_p_strobe_in_signal                                                                 => CONNECTED_TO_spwc_a_lvds_spw_lvds_p_strobe_in_signal,                                                                 --                                                                    .spw_lvds_p_strobe_in_signal
			spwc_a_lvds_spw_lvds_n_strobe_in_signal                                                                 => CONNECTED_TO_spwc_a_lvds_spw_lvds_n_strobe_in_signal,                                                                 --                                                                    .spw_lvds_n_strobe_in_signal
			spwc_b_enable_spw_rx_enable_signal                                                                      => CONNECTED_TO_spwc_b_enable_spw_rx_enable_signal,                                                                      --                                                       spwc_b_enable.spw_rx_enable_signal
			spwc_b_enable_spw_tx_enable_signal                                                                      => CONNECTED_TO_spwc_b_enable_spw_tx_enable_signal,                                                                      --                                                                    .spw_tx_enable_signal
			spwc_b_leds_spw_red_status_led_signal                                                                   => CONNECTED_TO_spwc_b_leds_spw_red_status_led_signal,                                                                   --                                                         spwc_b_leds.spw_red_status_led_signal
			spwc_b_leds_spw_green_status_led_signal                                                                 => CONNECTED_TO_spwc_b_leds_spw_green_status_led_signal,                                                                 --                                                                    .spw_green_status_led_signal
			spwc_b_lvds_spw_lvds_p_data_in_signal                                                                   => CONNECTED_TO_spwc_b_lvds_spw_lvds_p_data_in_signal,                                                                   --                                                         spwc_b_lvds.spw_lvds_p_data_in_signal
			spwc_b_lvds_spw_lvds_n_data_in_signal                                                                   => CONNECTED_TO_spwc_b_lvds_spw_lvds_n_data_in_signal,                                                                   --                                                                    .spw_lvds_n_data_in_signal
			spwc_b_lvds_spw_lvds_p_data_out_signal                                                                  => CONNECTED_TO_spwc_b_lvds_spw_lvds_p_data_out_signal,                                                                  --                                                                    .spw_lvds_p_data_out_signal
			spwc_b_lvds_spw_lvds_n_data_out_signal                                                                  => CONNECTED_TO_spwc_b_lvds_spw_lvds_n_data_out_signal,                                                                  --                                                                    .spw_lvds_n_data_out_signal
			spwc_b_lvds_spw_lvds_p_strobe_out_signal                                                                => CONNECTED_TO_spwc_b_lvds_spw_lvds_p_strobe_out_signal,                                                                --                                                                    .spw_lvds_p_strobe_out_signal
			spwc_b_lvds_spw_lvds_n_strobe_out_signal                                                                => CONNECTED_TO_spwc_b_lvds_spw_lvds_n_strobe_out_signal,                                                                --                                                                    .spw_lvds_n_strobe_out_signal
			spwc_b_lvds_spw_lvds_p_strobe_in_signal                                                                 => CONNECTED_TO_spwc_b_lvds_spw_lvds_p_strobe_in_signal,                                                                 --                                                                    .spw_lvds_p_strobe_in_signal
			spwc_b_lvds_spw_lvds_n_strobe_in_signal                                                                 => CONNECTED_TO_spwc_b_lvds_spw_lvds_n_strobe_in_signal,                                                                 --                                                                    .spw_lvds_n_strobe_in_signal
			spwc_c_enable_spw_rx_enable_signal                                                                      => CONNECTED_TO_spwc_c_enable_spw_rx_enable_signal,                                                                      --                                                       spwc_c_enable.spw_rx_enable_signal
			spwc_c_enable_spw_tx_enable_signal                                                                      => CONNECTED_TO_spwc_c_enable_spw_tx_enable_signal,                                                                      --                                                                    .spw_tx_enable_signal
			spwc_c_leds_spw_red_status_led_signal                                                                   => CONNECTED_TO_spwc_c_leds_spw_red_status_led_signal,                                                                   --                                                         spwc_c_leds.spw_red_status_led_signal
			spwc_c_leds_spw_green_status_led_signal                                                                 => CONNECTED_TO_spwc_c_leds_spw_green_status_led_signal,                                                                 --                                                                    .spw_green_status_led_signal
			spwc_c_lvds_spw_lvds_p_data_in_signal                                                                   => CONNECTED_TO_spwc_c_lvds_spw_lvds_p_data_in_signal,                                                                   --                                                         spwc_c_lvds.spw_lvds_p_data_in_signal
			spwc_c_lvds_spw_lvds_n_data_in_signal                                                                   => CONNECTED_TO_spwc_c_lvds_spw_lvds_n_data_in_signal,                                                                   --                                                                    .spw_lvds_n_data_in_signal
			spwc_c_lvds_spw_lvds_p_data_out_signal                                                                  => CONNECTED_TO_spwc_c_lvds_spw_lvds_p_data_out_signal,                                                                  --                                                                    .spw_lvds_p_data_out_signal
			spwc_c_lvds_spw_lvds_n_data_out_signal                                                                  => CONNECTED_TO_spwc_c_lvds_spw_lvds_n_data_out_signal,                                                                  --                                                                    .spw_lvds_n_data_out_signal
			spwc_c_lvds_spw_lvds_p_strobe_out_signal                                                                => CONNECTED_TO_spwc_c_lvds_spw_lvds_p_strobe_out_signal,                                                                --                                                                    .spw_lvds_p_strobe_out_signal
			spwc_c_lvds_spw_lvds_n_strobe_out_signal                                                                => CONNECTED_TO_spwc_c_lvds_spw_lvds_n_strobe_out_signal,                                                                --                                                                    .spw_lvds_n_strobe_out_signal
			spwc_c_lvds_spw_lvds_p_strobe_in_signal                                                                 => CONNECTED_TO_spwc_c_lvds_spw_lvds_p_strobe_in_signal,                                                                 --                                                                    .spw_lvds_p_strobe_in_signal
			spwc_c_lvds_spw_lvds_n_strobe_in_signal                                                                 => CONNECTED_TO_spwc_c_lvds_spw_lvds_n_strobe_in_signal,                                                                 --                                                                    .spw_lvds_n_strobe_in_signal
			spwc_d_enable_spw_rx_enable_signal                                                                      => CONNECTED_TO_spwc_d_enable_spw_rx_enable_signal,                                                                      --                                                       spwc_d_enable.spw_rx_enable_signal
			spwc_d_enable_spw_tx_enable_signal                                                                      => CONNECTED_TO_spwc_d_enable_spw_tx_enable_signal,                                                                      --                                                                    .spw_tx_enable_signal
			spwc_d_leds_spw_red_status_led_signal                                                                   => CONNECTED_TO_spwc_d_leds_spw_red_status_led_signal,                                                                   --                                                         spwc_d_leds.spw_red_status_led_signal
			spwc_d_leds_spw_green_status_led_signal                                                                 => CONNECTED_TO_spwc_d_leds_spw_green_status_led_signal,                                                                 --                                                                    .spw_green_status_led_signal
			spwc_d_lvds_spw_lvds_p_data_in_signal                                                                   => CONNECTED_TO_spwc_d_lvds_spw_lvds_p_data_in_signal,                                                                   --                                                         spwc_d_lvds.spw_lvds_p_data_in_signal
			spwc_d_lvds_spw_lvds_n_data_in_signal                                                                   => CONNECTED_TO_spwc_d_lvds_spw_lvds_n_data_in_signal,                                                                   --                                                                    .spw_lvds_n_data_in_signal
			spwc_d_lvds_spw_lvds_p_data_out_signal                                                                  => CONNECTED_TO_spwc_d_lvds_spw_lvds_p_data_out_signal,                                                                  --                                                                    .spw_lvds_p_data_out_signal
			spwc_d_lvds_spw_lvds_n_data_out_signal                                                                  => CONNECTED_TO_spwc_d_lvds_spw_lvds_n_data_out_signal,                                                                  --                                                                    .spw_lvds_n_data_out_signal
			spwc_d_lvds_spw_lvds_p_strobe_out_signal                                                                => CONNECTED_TO_spwc_d_lvds_spw_lvds_p_strobe_out_signal,                                                                --                                                                    .spw_lvds_p_strobe_out_signal
			spwc_d_lvds_spw_lvds_n_strobe_out_signal                                                                => CONNECTED_TO_spwc_d_lvds_spw_lvds_n_strobe_out_signal,                                                                --                                                                    .spw_lvds_n_strobe_out_signal
			spwc_d_lvds_spw_lvds_p_strobe_in_signal                                                                 => CONNECTED_TO_spwc_d_lvds_spw_lvds_p_strobe_in_signal,                                                                 --                                                                    .spw_lvds_p_strobe_in_signal
			spwc_d_lvds_spw_lvds_n_strobe_in_signal                                                                 => CONNECTED_TO_spwc_d_lvds_spw_lvds_n_strobe_in_signal,                                                                 --                                                                    .spw_lvds_n_strobe_in_signal
			spwc_e_enable_spw_rx_enable_signal                                                                      => CONNECTED_TO_spwc_e_enable_spw_rx_enable_signal,                                                                      --                                                       spwc_e_enable.spw_rx_enable_signal
			spwc_e_enable_spw_tx_enable_signal                                                                      => CONNECTED_TO_spwc_e_enable_spw_tx_enable_signal,                                                                      --                                                                    .spw_tx_enable_signal
			spwc_e_leds_spw_red_status_led_signal                                                                   => CONNECTED_TO_spwc_e_leds_spw_red_status_led_signal,                                                                   --                                                         spwc_e_leds.spw_red_status_led_signal
			spwc_e_leds_spw_green_status_led_signal                                                                 => CONNECTED_TO_spwc_e_leds_spw_green_status_led_signal,                                                                 --                                                                    .spw_green_status_led_signal
			spwc_e_lvds_spw_lvds_p_data_in_signal                                                                   => CONNECTED_TO_spwc_e_lvds_spw_lvds_p_data_in_signal,                                                                   --                                                         spwc_e_lvds.spw_lvds_p_data_in_signal
			spwc_e_lvds_spw_lvds_n_data_in_signal                                                                   => CONNECTED_TO_spwc_e_lvds_spw_lvds_n_data_in_signal,                                                                   --                                                                    .spw_lvds_n_data_in_signal
			spwc_e_lvds_spw_lvds_p_data_out_signal                                                                  => CONNECTED_TO_spwc_e_lvds_spw_lvds_p_data_out_signal,                                                                  --                                                                    .spw_lvds_p_data_out_signal
			spwc_e_lvds_spw_lvds_n_data_out_signal                                                                  => CONNECTED_TO_spwc_e_lvds_spw_lvds_n_data_out_signal,                                                                  --                                                                    .spw_lvds_n_data_out_signal
			spwc_e_lvds_spw_lvds_p_strobe_out_signal                                                                => CONNECTED_TO_spwc_e_lvds_spw_lvds_p_strobe_out_signal,                                                                --                                                                    .spw_lvds_p_strobe_out_signal
			spwc_e_lvds_spw_lvds_n_strobe_out_signal                                                                => CONNECTED_TO_spwc_e_lvds_spw_lvds_n_strobe_out_signal,                                                                --                                                                    .spw_lvds_n_strobe_out_signal
			spwc_e_lvds_spw_lvds_p_strobe_in_signal                                                                 => CONNECTED_TO_spwc_e_lvds_spw_lvds_p_strobe_in_signal,                                                                 --                                                                    .spw_lvds_p_strobe_in_signal
			spwc_e_lvds_spw_lvds_n_strobe_in_signal                                                                 => CONNECTED_TO_spwc_e_lvds_spw_lvds_n_strobe_in_signal,                                                                 --                                                                    .spw_lvds_n_strobe_in_signal
			spwc_f_enable_spw_rx_enable_signal                                                                      => CONNECTED_TO_spwc_f_enable_spw_rx_enable_signal,                                                                      --                                                       spwc_f_enable.spw_rx_enable_signal
			spwc_f_enable_spw_tx_enable_signal                                                                      => CONNECTED_TO_spwc_f_enable_spw_tx_enable_signal,                                                                      --                                                                    .spw_tx_enable_signal
			spwc_f_leds_spw_red_status_led_signal                                                                   => CONNECTED_TO_spwc_f_leds_spw_red_status_led_signal,                                                                   --                                                         spwc_f_leds.spw_red_status_led_signal
			spwc_f_leds_spw_green_status_led_signal                                                                 => CONNECTED_TO_spwc_f_leds_spw_green_status_led_signal,                                                                 --                                                                    .spw_green_status_led_signal
			spwc_f_lvds_spw_lvds_p_data_in_signal                                                                   => CONNECTED_TO_spwc_f_lvds_spw_lvds_p_data_in_signal,                                                                   --                                                         spwc_f_lvds.spw_lvds_p_data_in_signal
			spwc_f_lvds_spw_lvds_n_data_in_signal                                                                   => CONNECTED_TO_spwc_f_lvds_spw_lvds_n_data_in_signal,                                                                   --                                                                    .spw_lvds_n_data_in_signal
			spwc_f_lvds_spw_lvds_p_data_out_signal                                                                  => CONNECTED_TO_spwc_f_lvds_spw_lvds_p_data_out_signal,                                                                  --                                                                    .spw_lvds_p_data_out_signal
			spwc_f_lvds_spw_lvds_n_data_out_signal                                                                  => CONNECTED_TO_spwc_f_lvds_spw_lvds_n_data_out_signal,                                                                  --                                                                    .spw_lvds_n_data_out_signal
			spwc_f_lvds_spw_lvds_p_strobe_out_signal                                                                => CONNECTED_TO_spwc_f_lvds_spw_lvds_p_strobe_out_signal,                                                                --                                                                    .spw_lvds_p_strobe_out_signal
			spwc_f_lvds_spw_lvds_n_strobe_out_signal                                                                => CONNECTED_TO_spwc_f_lvds_spw_lvds_n_strobe_out_signal,                                                                --                                                                    .spw_lvds_n_strobe_out_signal
			spwc_f_lvds_spw_lvds_p_strobe_in_signal                                                                 => CONNECTED_TO_spwc_f_lvds_spw_lvds_p_strobe_in_signal,                                                                 --                                                                    .spw_lvds_p_strobe_in_signal
			spwc_f_lvds_spw_lvds_n_strobe_in_signal                                                                 => CONNECTED_TO_spwc_f_lvds_spw_lvds_n_strobe_in_signal,                                                                 --                                                                    .spw_lvds_n_strobe_in_signal
			spwc_g_enable_spw_rx_enable_signal                                                                      => CONNECTED_TO_spwc_g_enable_spw_rx_enable_signal,                                                                      --                                                       spwc_g_enable.spw_rx_enable_signal
			spwc_g_enable_spw_tx_enable_signal                                                                      => CONNECTED_TO_spwc_g_enable_spw_tx_enable_signal,                                                                      --                                                                    .spw_tx_enable_signal
			spwc_g_leds_spw_red_status_led_signal                                                                   => CONNECTED_TO_spwc_g_leds_spw_red_status_led_signal,                                                                   --                                                         spwc_g_leds.spw_red_status_led_signal
			spwc_g_leds_spw_green_status_led_signal                                                                 => CONNECTED_TO_spwc_g_leds_spw_green_status_led_signal,                                                                 --                                                                    .spw_green_status_led_signal
			spwc_g_lvds_spw_lvds_p_data_in_signal                                                                   => CONNECTED_TO_spwc_g_lvds_spw_lvds_p_data_in_signal,                                                                   --                                                         spwc_g_lvds.spw_lvds_p_data_in_signal
			spwc_g_lvds_spw_lvds_n_data_in_signal                                                                   => CONNECTED_TO_spwc_g_lvds_spw_lvds_n_data_in_signal,                                                                   --                                                                    .spw_lvds_n_data_in_signal
			spwc_g_lvds_spw_lvds_p_data_out_signal                                                                  => CONNECTED_TO_spwc_g_lvds_spw_lvds_p_data_out_signal,                                                                  --                                                                    .spw_lvds_p_data_out_signal
			spwc_g_lvds_spw_lvds_n_data_out_signal                                                                  => CONNECTED_TO_spwc_g_lvds_spw_lvds_n_data_out_signal,                                                                  --                                                                    .spw_lvds_n_data_out_signal
			spwc_g_lvds_spw_lvds_p_strobe_out_signal                                                                => CONNECTED_TO_spwc_g_lvds_spw_lvds_p_strobe_out_signal,                                                                --                                                                    .spw_lvds_p_strobe_out_signal
			spwc_g_lvds_spw_lvds_n_strobe_out_signal                                                                => CONNECTED_TO_spwc_g_lvds_spw_lvds_n_strobe_out_signal,                                                                --                                                                    .spw_lvds_n_strobe_out_signal
			spwc_g_lvds_spw_lvds_p_strobe_in_signal                                                                 => CONNECTED_TO_spwc_g_lvds_spw_lvds_p_strobe_in_signal,                                                                 --                                                                    .spw_lvds_p_strobe_in_signal
			spwc_g_lvds_spw_lvds_n_strobe_in_signal                                                                 => CONNECTED_TO_spwc_g_lvds_spw_lvds_n_strobe_in_signal,                                                                 --                                                                    .spw_lvds_n_strobe_in_signal
			spwc_h_enable_spw_rx_enable_signal                                                                      => CONNECTED_TO_spwc_h_enable_spw_rx_enable_signal,                                                                      --                                                       spwc_h_enable.spw_rx_enable_signal
			spwc_h_enable_spw_tx_enable_signal                                                                      => CONNECTED_TO_spwc_h_enable_spw_tx_enable_signal,                                                                      --                                                                    .spw_tx_enable_signal
			spwc_h_leds_spw_red_status_led_signal                                                                   => CONNECTED_TO_spwc_h_leds_spw_red_status_led_signal,                                                                   --                                                         spwc_h_leds.spw_red_status_led_signal
			spwc_h_leds_spw_green_status_led_signal                                                                 => CONNECTED_TO_spwc_h_leds_spw_green_status_led_signal,                                                                 --                                                                    .spw_green_status_led_signal
			spwc_h_lvds_spw_lvds_p_data_in_signal                                                                   => CONNECTED_TO_spwc_h_lvds_spw_lvds_p_data_in_signal,                                                                   --                                                         spwc_h_lvds.spw_lvds_p_data_in_signal
			spwc_h_lvds_spw_lvds_n_data_in_signal                                                                   => CONNECTED_TO_spwc_h_lvds_spw_lvds_n_data_in_signal,                                                                   --                                                                    .spw_lvds_n_data_in_signal
			spwc_h_lvds_spw_lvds_p_data_out_signal                                                                  => CONNECTED_TO_spwc_h_lvds_spw_lvds_p_data_out_signal,                                                                  --                                                                    .spw_lvds_p_data_out_signal
			spwc_h_lvds_spw_lvds_n_data_out_signal                                                                  => CONNECTED_TO_spwc_h_lvds_spw_lvds_n_data_out_signal,                                                                  --                                                                    .spw_lvds_n_data_out_signal
			spwc_h_lvds_spw_lvds_p_strobe_out_signal                                                                => CONNECTED_TO_spwc_h_lvds_spw_lvds_p_strobe_out_signal,                                                                --                                                                    .spw_lvds_p_strobe_out_signal
			spwc_h_lvds_spw_lvds_n_strobe_out_signal                                                                => CONNECTED_TO_spwc_h_lvds_spw_lvds_n_strobe_out_signal,                                                                --                                                                    .spw_lvds_n_strobe_out_signal
			spwc_h_lvds_spw_lvds_p_strobe_in_signal                                                                 => CONNECTED_TO_spwc_h_lvds_spw_lvds_p_strobe_in_signal,                                                                 --                                                                    .spw_lvds_p_strobe_in_signal
			spwc_h_lvds_spw_lvds_n_strobe_in_signal                                                                 => CONNECTED_TO_spwc_h_lvds_spw_lvds_n_strobe_in_signal,                                                                 --                                                                    .spw_lvds_n_strobe_in_signal
			spwm_h_select_mux_select_signal                                                                         => CONNECTED_TO_spwm_h_select_mux_select_signal,                                                                         --                                                       spwm_h_select.mux_select_signal
			ssdp_ssdp0                                                                                              => CONNECTED_TO_ssdp_ssdp0,                                                                                              --                                                                ssdp.ssdp0
			ssdp_ssdp1                                                                                              => CONNECTED_TO_ssdp_ssdp1,                                                                                              --                                                                    .ssdp1
			sync_in_conduit                                                                                         => CONNECTED_TO_sync_in_conduit,                                                                                         --                                                             sync_in.conduit
			sync_in_en_conduit                                                                                      => CONNECTED_TO_sync_in_en_conduit,                                                                                      --                                                          sync_in_en.conduit
			sync_out_conduit                                                                                        => CONNECTED_TO_sync_out_conduit,                                                                                        --                                                            sync_out.conduit
			sync_out_en_conduit                                                                                     => CONNECTED_TO_sync_out_en_conduit,                                                                                     --                                                         sync_out_en.conduit
			sync_spw1_conduit                                                                                       => CONNECTED_TO_sync_spw1_conduit,                                                                                       --                                                           sync_spw1.conduit
			sync_spw2_conduit                                                                                       => CONNECTED_TO_sync_spw2_conduit,                                                                                       --                                                           sync_spw2.conduit
			sync_spw3_conduit                                                                                       => CONNECTED_TO_sync_spw3_conduit,                                                                                       --                                                           sync_spw3.conduit
			sync_spw4_conduit                                                                                       => CONNECTED_TO_sync_spw4_conduit,                                                                                       --                                                           sync_spw4.conduit
			sync_spw5_conduit                                                                                       => CONNECTED_TO_sync_spw5_conduit,                                                                                       --                                                           sync_spw5.conduit
			sync_spw6_conduit                                                                                       => CONNECTED_TO_sync_spw6_conduit,                                                                                       --                                                           sync_spw6.conduit
			sync_spw7_conduit                                                                                       => CONNECTED_TO_sync_spw7_conduit,                                                                                       --                                                           sync_spw7.conduit
			sync_spw8_conduit                                                                                       => CONNECTED_TO_sync_spw8_conduit,                                                                                       --                                                           sync_spw8.conduit
			temp_scl_export                                                                                         => CONNECTED_TO_temp_scl_export,                                                                                         --                                                            temp_scl.export
			temp_sda_export                                                                                         => CONNECTED_TO_temp_sda_export,                                                                                         --                                                            temp_sda.export
			timer_1ms_external_port_export                                                                          => CONNECTED_TO_timer_1ms_external_port_export,                                                                          --                                             timer_1ms_external_port.export
			timer_1us_external_port_export                                                                          => CONNECTED_TO_timer_1us_external_port_export,                                                                          --                                             timer_1us_external_port.export
			tristate_conduit_tcm_address_out                                                                        => CONNECTED_TO_tristate_conduit_tcm_address_out,                                                                        --                                                    tristate_conduit.tcm_address_out
			tristate_conduit_tcm_read_n_out                                                                         => CONNECTED_TO_tristate_conduit_tcm_read_n_out,                                                                         --                                                                    .tcm_read_n_out
			tristate_conduit_tcm_write_n_out                                                                        => CONNECTED_TO_tristate_conduit_tcm_write_n_out,                                                                        --                                                                    .tcm_write_n_out
			tristate_conduit_tcm_data_out                                                                           => CONNECTED_TO_tristate_conduit_tcm_data_out,                                                                           --                                                                    .tcm_data_out
			tristate_conduit_tcm_chipselect_n_out                                                                   => CONNECTED_TO_tristate_conduit_tcm_chipselect_n_out,                                                                   --                                                                    .tcm_chipselect_n_out
			umft601a_pins_umft_clock_signal                                                                         => CONNECTED_TO_umft601a_pins_umft_clock_signal,                                                                         --                                                       umft601a_pins.umft_clock_signal
			umft601a_pins_umft_txe_n_signal                                                                         => CONNECTED_TO_umft601a_pins_umft_txe_n_signal,                                                                         --                                                                    .umft_txe_n_signal
			umft601a_pins_umft_rxf_n_signal                                                                         => CONNECTED_TO_umft601a_pins_umft_rxf_n_signal,                                                                         --                                                                    .umft_rxf_n_signal
			umft601a_pins_umft_data_signal                                                                          => CONNECTED_TO_umft601a_pins_umft_data_signal,                                                                          --                                                                    .umft_data_signal
			umft601a_pins_umft_be_signal                                                                            => CONNECTED_TO_umft601a_pins_umft_be_signal,                                                                            --                                                                    .umft_be_signal
			umft601a_pins_umft_wakeup_n_signal                                                                      => CONNECTED_TO_umft601a_pins_umft_wakeup_n_signal,                                                                      --                                                                    .umft_wakeup_n_signal
			umft601a_pins_umft_gpio_bus_signal                                                                      => CONNECTED_TO_umft601a_pins_umft_gpio_bus_signal,                                                                      --                                                                    .umft_gpio_bus_signal
			umft601a_pins_umft_reset_n_signal                                                                       => CONNECTED_TO_umft601a_pins_umft_reset_n_signal,                                                                       --                                                                    .umft_reset_n_signal
			umft601a_pins_umft_wr_n_signal                                                                          => CONNECTED_TO_umft601a_pins_umft_wr_n_signal,                                                                          --                                                                    .umft_wr_n_signal
			umft601a_pins_umft_rd_n_signal                                                                          => CONNECTED_TO_umft601a_pins_umft_rd_n_signal,                                                                          --                                                                    .umft_rd_n_signal
			umft601a_pins_umft_oe_n_signal                                                                          => CONNECTED_TO_umft601a_pins_umft_oe_n_signal,                                                                          --                                                                    .umft_oe_n_signal
			umft601a_pins_umft_siwu_n_signal                                                                        => CONNECTED_TO_umft601a_pins_umft_siwu_n_signal                                                                         --                                                                    .umft_siwu_n_signal
		);

