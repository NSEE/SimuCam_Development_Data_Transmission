library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity avalon_mm_data_buffer_write_ent is
	port(
		clk : in std_logic;
		rst : in std_logic
	);
end entity avalon_mm_data_buffer_write_ent;

architecture RTL of avalon_mm_data_buffer_write_ent is
	
begin

end architecture RTL;
