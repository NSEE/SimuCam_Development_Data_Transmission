package data_buffer_pkg is
	
end package data_buffer_pkg;

package body data_buffer_pkg is
	
end package body data_buffer_pkg;
