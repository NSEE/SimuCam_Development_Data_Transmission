-- MebX_Qsys_Project.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity MebX_Qsys_Project is
	port (
		clk50_clk                                  : in  std_logic                     := '0';             --                          clk50.clk
		rs232_uart_rxd                             : in  std_logic                     := '0';             --                     rs232_uart.rxd
		rs232_uart_txd                             : out std_logic;                                        --                               .txd
		rs232_uart_cts_n                           : in  std_logic                     := '0';             --                               .cts_n
		rs232_uart_rts_n                           : out std_logic;                                        --                               .rts_n
		rs232_uart_irq_irq                         : out std_logic;                                        --                 rs232_uart_irq.irq
		rst_reset_n                                : in  std_logic                     := '0';             --                            rst.reset_n
		uart_module_uart_txd_signal                : out std_logic;                                        --                    uart_module.uart_txd_signal
		uart_module_uart_rxd_signal                : in  std_logic                     := '0';             --                               .uart_rxd_signal
		uart_module_uart_rts_signal                : in  std_logic                     := '0';             --                               .uart_rts_signal
		uart_module_uart_cts_signal                : out std_logic;                                        --                               .uart_cts_signal
		uart_module_top_0_avalon_slave_address     : in  std_logic_vector(7 downto 0)  := (others => '0'); -- uart_module_top_0_avalon_slave.address
		uart_module_top_0_avalon_slave_read        : in  std_logic                     := '0';             --                               .read
		uart_module_top_0_avalon_slave_write       : in  std_logic                     := '0';             --                               .write
		uart_module_top_0_avalon_slave_waitrequest : out std_logic;                                        --                               .waitrequest
		uart_module_top_0_avalon_slave_writedata   : in  std_logic_vector(31 downto 0) := (others => '0'); --                               .writedata
		uart_module_top_0_avalon_slave_readdata    : out std_logic_vector(31 downto 0)                     --                               .readdata
	);
end entity MebX_Qsys_Project;

architecture rtl of MebX_Qsys_Project is
	component MebX_Qsys_Project_rs232_uart is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			cts_n         : in  std_logic                     := 'X';             -- export
			rts_n         : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component MebX_Qsys_Project_rs232_uart;

	component uart_module_top is
		port (
			reset_sink_reset          : in  std_logic                     := 'X';             -- reset
			clock_sink_clk            : in  std_logic                     := 'X';             -- clk
			uart_txd                  : out std_logic;                                        -- uart_txd_signal
			uart_rxd                  : in  std_logic                     := 'X';             -- uart_rxd_signal
			uart_rts                  : in  std_logic                     := 'X';             -- uart_rts_signal
			uart_cts                  : out std_logic;                                        -- uart_cts_signal
			avalon_slave_address      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			avalon_slave_read         : in  std_logic                     := 'X';             -- read
			avalon_slave_write        : in  std_logic                     := 'X';             -- write
			avalon_slave_waitrequest  : out std_logic;                                        -- waitrequest
			avalon_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalon_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			avalon_master_address     : out std_logic_vector(5 downto 0);                     -- address
			avalon_master_read        : out std_logic;                                        -- read
			avalon_master_write       : out std_logic;                                        -- write
			avalon_master_writedata   : out std_logic_vector(15 downto 0);                    -- writedata
			avalon_master_readdata    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			avalon_master_waitrequest : in  std_logic                     := 'X'              -- waitrequest
		);
	end component uart_module_top;

	component MebX_Qsys_Project_mm_interconnect_0 is
		port (
			clk_50_clk_clk                                           : in  std_logic                     := 'X';             -- clk
			uart_module_top_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			uart_module_top_0_avalon_master_address                  : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			uart_module_top_0_avalon_master_waitrequest              : out std_logic;                                        -- waitrequest
			uart_module_top_0_avalon_master_read                     : in  std_logic                     := 'X';             -- read
			uart_module_top_0_avalon_master_readdata                 : out std_logic_vector(15 downto 0);                    -- readdata
			uart_module_top_0_avalon_master_write                    : in  std_logic                     := 'X';             -- write
			uart_module_top_0_avalon_master_writedata                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			rs232_uart_s1_address                                    : out std_logic_vector(2 downto 0);                     -- address
			rs232_uart_s1_write                                      : out std_logic;                                        -- write
			rs232_uart_s1_read                                       : out std_logic;                                        -- read
			rs232_uart_s1_readdata                                   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			rs232_uart_s1_writedata                                  : out std_logic_vector(15 downto 0);                    -- writedata
			rs232_uart_s1_begintransfer                              : out std_logic;                                        -- begintransfer
			rs232_uart_s1_chipselect                                 : out std_logic                                         -- chipselect
		);
	end component MebX_Qsys_Project_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal uart_module_top_0_avalon_master_readdata        : std_logic_vector(15 downto 0); -- mm_interconnect_0:uart_module_top_0_avalon_master_readdata -> uart_module_top_0:avalon_master_readdata
	signal uart_module_top_0_avalon_master_waitrequest     : std_logic;                     -- mm_interconnect_0:uart_module_top_0_avalon_master_waitrequest -> uart_module_top_0:avalon_master_waitrequest
	signal uart_module_top_0_avalon_master_address         : std_logic_vector(5 downto 0);  -- uart_module_top_0:avalon_master_address -> mm_interconnect_0:uart_module_top_0_avalon_master_address
	signal uart_module_top_0_avalon_master_read            : std_logic;                     -- uart_module_top_0:avalon_master_read -> mm_interconnect_0:uart_module_top_0_avalon_master_read
	signal uart_module_top_0_avalon_master_write           : std_logic;                     -- uart_module_top_0:avalon_master_write -> mm_interconnect_0:uart_module_top_0_avalon_master_write
	signal uart_module_top_0_avalon_master_writedata       : std_logic_vector(15 downto 0); -- uart_module_top_0:avalon_master_writedata -> mm_interconnect_0:uart_module_top_0_avalon_master_writedata
	signal mm_interconnect_0_rs232_uart_s1_chipselect      : std_logic;                     -- mm_interconnect_0:rs232_uart_s1_chipselect -> rs232_uart:chipselect
	signal mm_interconnect_0_rs232_uart_s1_readdata        : std_logic_vector(15 downto 0); -- rs232_uart:readdata -> mm_interconnect_0:rs232_uart_s1_readdata
	signal mm_interconnect_0_rs232_uart_s1_address         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:rs232_uart_s1_address -> rs232_uart:address
	signal mm_interconnect_0_rs232_uart_s1_read            : std_logic;                     -- mm_interconnect_0:rs232_uart_s1_read -> mm_interconnect_0_rs232_uart_s1_read:in
	signal mm_interconnect_0_rs232_uart_s1_begintransfer   : std_logic;                     -- mm_interconnect_0:rs232_uart_s1_begintransfer -> rs232_uart:begintransfer
	signal mm_interconnect_0_rs232_uart_s1_write           : std_logic;                     -- mm_interconnect_0:rs232_uart_s1_write -> mm_interconnect_0_rs232_uart_s1_write:in
	signal mm_interconnect_0_rs232_uart_s1_writedata       : std_logic_vector(15 downto 0); -- mm_interconnect_0:rs232_uart_s1_writedata -> rs232_uart:writedata
	signal rst_controller_reset_out_reset                  : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:uart_module_top_0_reset_sink_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, uart_module_top_0:reset_sink_reset]
	signal rst_reset_n_ports_inv                           : std_logic;                     -- rst_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_rs232_uart_s1_read_ports_inv  : std_logic;                     -- mm_interconnect_0_rs232_uart_s1_read:inv -> rs232_uart:read_n
	signal mm_interconnect_0_rs232_uart_s1_write_ports_inv : std_logic;                     -- mm_interconnect_0_rs232_uart_s1_write:inv -> rs232_uart:write_n
	signal rst_controller_reset_out_reset_ports_inv        : std_logic;                     -- rst_controller_reset_out_reset:inv -> rs232_uart:reset_n

begin

	rs232_uart : component MebX_Qsys_Project_rs232_uart
		port map (
			clk           => clk50_clk,                                       --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address       => mm_interconnect_0_rs232_uart_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_rs232_uart_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_rs232_uart_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_rs232_uart_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_rs232_uart_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_rs232_uart_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_rs232_uart_s1_readdata,        --                    .readdata
			rxd           => rs232_uart_rxd,                                  -- external_connection.export
			txd           => rs232_uart_txd,                                  --                    .export
			cts_n         => rs232_uart_cts_n,                                --                    .export
			rts_n         => rs232_uart_rts_n,                                --                    .export
			irq           => rs232_uart_irq_irq                               --                 irq.irq
		);

	uart_module_top_0 : component uart_module_top
		port map (
			reset_sink_reset          => rst_controller_reset_out_reset,              --    reset_sink.reset
			clock_sink_clk            => clk50_clk,                                   --    clock_sink.clk
			uart_txd                  => uart_module_uart_txd_signal,                 --   conduit_end.uart_txd_signal
			uart_rxd                  => uart_module_uart_rxd_signal,                 --              .uart_rxd_signal
			uart_rts                  => uart_module_uart_rts_signal,                 --              .uart_rts_signal
			uart_cts                  => uart_module_uart_cts_signal,                 --              .uart_cts_signal
			avalon_slave_address      => uart_module_top_0_avalon_slave_address,      --  avalon_slave.address
			avalon_slave_read         => uart_module_top_0_avalon_slave_read,         --              .read
			avalon_slave_write        => uart_module_top_0_avalon_slave_write,        --              .write
			avalon_slave_waitrequest  => uart_module_top_0_avalon_slave_waitrequest,  --              .waitrequest
			avalon_slave_writedata    => uart_module_top_0_avalon_slave_writedata,    --              .writedata
			avalon_slave_readdata     => uart_module_top_0_avalon_slave_readdata,     --              .readdata
			avalon_master_address     => uart_module_top_0_avalon_master_address,     -- avalon_master.address
			avalon_master_read        => uart_module_top_0_avalon_master_read,        --              .read
			avalon_master_write       => uart_module_top_0_avalon_master_write,       --              .write
			avalon_master_writedata   => uart_module_top_0_avalon_master_writedata,   --              .writedata
			avalon_master_readdata    => uart_module_top_0_avalon_master_readdata,    --              .readdata
			avalon_master_waitrequest => uart_module_top_0_avalon_master_waitrequest  --              .waitrequest
		);

	mm_interconnect_0 : component MebX_Qsys_Project_mm_interconnect_0
		port map (
			clk_50_clk_clk                                           => clk50_clk,                                     --                                         clk_50_clk.clk
			uart_module_top_0_reset_sink_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                -- uart_module_top_0_reset_sink_reset_bridge_in_reset.reset
			uart_module_top_0_avalon_master_address                  => uart_module_top_0_avalon_master_address,       --                    uart_module_top_0_avalon_master.address
			uart_module_top_0_avalon_master_waitrequest              => uart_module_top_0_avalon_master_waitrequest,   --                                                   .waitrequest
			uart_module_top_0_avalon_master_read                     => uart_module_top_0_avalon_master_read,          --                                                   .read
			uart_module_top_0_avalon_master_readdata                 => uart_module_top_0_avalon_master_readdata,      --                                                   .readdata
			uart_module_top_0_avalon_master_write                    => uart_module_top_0_avalon_master_write,         --                                                   .write
			uart_module_top_0_avalon_master_writedata                => uart_module_top_0_avalon_master_writedata,     --                                                   .writedata
			rs232_uart_s1_address                                    => mm_interconnect_0_rs232_uart_s1_address,       --                                      rs232_uart_s1.address
			rs232_uart_s1_write                                      => mm_interconnect_0_rs232_uart_s1_write,         --                                                   .write
			rs232_uart_s1_read                                       => mm_interconnect_0_rs232_uart_s1_read,          --                                                   .read
			rs232_uart_s1_readdata                                   => mm_interconnect_0_rs232_uart_s1_readdata,      --                                                   .readdata
			rs232_uart_s1_writedata                                  => mm_interconnect_0_rs232_uart_s1_writedata,     --                                                   .writedata
			rs232_uart_s1_begintransfer                              => mm_interconnect_0_rs232_uart_s1_begintransfer, --                                                   .begintransfer
			rs232_uart_s1_chipselect                                 => mm_interconnect_0_rs232_uart_s1_chipselect     --                                                   .chipselect
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,          -- reset_in0.reset
			clk            => clk50_clk,                      --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_reset_n_ports_inv <= not rst_reset_n;

	mm_interconnect_0_rs232_uart_s1_read_ports_inv <= not mm_interconnect_0_rs232_uart_s1_read;

	mm_interconnect_0_rs232_uart_s1_write_ports_inv <= not mm_interconnect_0_rs232_uart_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of MebX_Qsys_Project
