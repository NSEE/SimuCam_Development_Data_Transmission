package data_controller_pkg is
	
end package data_controller_pkg;

package body data_controller_pkg is
	
end package body data_controller_pkg;
