library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity data_scheduler_ent is
	port(
		clk_i : in std_logic;
		rst_i : in std_logic
	);
end entity data_scheduler_ent;

architecture RTL of data_scheduler_ent is
	
begin

end architecture RTL;
