package data_scheduler_pkg is
	
end package data_scheduler_pkg;

package body data_scheduler_pkg is
	
end package body data_scheduler_pkg;
