// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:49 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cJfRo8+eqRm3g0WImZivAiVuXErQBdkQJ1DNh/2wft8QMiAbQyaufG0lHW1kqavm
BjcWduhP7481N0Ar+2wCM12D70y/aQI61dkwUDtYZhOym5R8NaWHJUkTxG+q/shP
amTZivc2d3Bi6Xy0tA1tBwpPlIGJZo/8BobzYXTArrc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21712)
hR90Fd9fpXn/PwVLf4wFSpkwYbd9+/jOrKLBq5zERgqbbX57IfUHY/pLGuPKaEf6
mVXIMiu1P3zdnCyNgr2khnrZ7fOzGwHjuuu475R9RIxJtF1nfA15xw5OyKJ//WXd
/2Ft2YL1/ZUwAFFgPftBS2lwFPJ8d3NV8eVRbKMypqWct1VTXCVPDWz3vdpcgITr
PSSfiLwfc8Z89XhU7OgyJYMvsemk3sV1zQNjkztxedMHo9UHPqXOKrdYUPfdJy99
vE+mxd56sV5dA8MTO+w3h1Jj3QmUMQnXYzYlMf2jb/yCil+XWpQuT/Lb9Ch73MA3
3M8KEjaLvBlPjKVdimIm7/NYwW6aiEoAwjWwEkq3/yzys1uumQrvsbVDyKRskT8O
wT7mfAdbOrXIeS8w1TNR54SDMqETXd1xmtuatNSyP79XORpkfVUdA1VjdBhMlP0m
BLElYYPPE/7yZudgCBl7zyQV5QRbrnXvat2vVLTZZ8I7NQ1AXjXP6m2TA94t928m
exomvrgjBjrz8Mf6vcU+hmILj+SAGNuXKofcBMHQWqogWa9w8Oq9B4s1h9V4sWBy
ARE22d01JwX9gN3iTaA825FW76Kr3ax2YkPmrOT7qfblzEgEjy8qlbMap56NJ+l6
qWg8NWS3d13YbwSpes2m2iG5FMMYKwGNm0nus/fAHF+BiCTcO5JI5OOfXWqjc7+V
vUdK8tKdUR+4xkQvsOD1dbSIhOh8leJ3BM9KKjayLBBe7fCEL0cK1PuvgdzFilCL
UluxqWLfzczjYioyqdidp3kDzGvlGP7TZdWG0HAuR8kt+EWMQ0Q/8Zi6b+nJNC85
r/T8LwbLYLIWyK60Ew0iiC6I134gebJZZ2lyByHEqibHEkaYULNkj+GtxR3SM4Xq
y+QOtJgISjJVfLywrXGztVdRpi2vxNdkba87clyQv5tPKLvLyf9QnEUF3/F8Q0kw
quhsG0otGW6p1HIe0F+CfK5kK2kdYFzst6USO13jwS7J+nePlMJV13wwYvEkGCb9
DRdNaAsFjt8ZRldSiS5/YgqoZzEcCvPuVd6SbPHLxjRCrfn7w7KSdbu/T7JbrcSb
Tmxm6f4mT7XVw42EL/PIzjRqgaWwSAh5U3wiFBsvNTmzhCQQLbyrF3zuhW3bKcyy
k3WzSWciDrWjWpSlgj4R8b8qMBwWZhwA4xeo1WcoORgXQ65SGSA8R424qbB8uLVB
kwhHR8DmTDTWFQzzjPtrQWx8guDi1szQ0I9tKYKuijB+mZ75Tj6UsZuB2LVSYrLx
tWIgQScyQYut0Jp/E3bgslFToNwRlPO+LxpthkvldkBxMU9GtU7/b4Yqg7pNH01A
2GQWAUl94TXzyrfALnqf+z96CmyFO98CWRs92cL8DULAgW+Zn9PIJtzTvY29Egrg
x2WChdoLQxAF2PyIWhSQJlbmKdTN9Srme4mKzVupcBDiu6Te85/50c96W1Lcabol
r8pkR1fjy/bR0w+PCPH3VUvau9ggcuaPcUbK6XOl18mBi8EJ9rV56R7Fn9onJreR
ZLRZ0WirwdZ+0QHkZAryThCa00tnIb9IpPdT2boo01zVhOrSJq58MISG/qD9p78q
w8u6x+sDw5n8JzOoKS9BkUQJKWMibq4I+TwL6yOm12XJHD8avDeqCog/yTr8i/Ht
oT+iD2CCq5LjS2bkpKXrvO/NvBPalHHDZoX1B5az+Ih+RjAaBAFfsTqCHBALWD1m
iC22Zp5cDnMONwX+l0RGrW6nPHraN4DJ99IkPqMTQWhfGiEiluBJkJ9U9hyi6vSN
Yf/9sjeCJXlbI8nUt+n3KbKm12DsS7+RcSYesVsR4K2k72zJVQDyhStkzh4GkO07
tivDNv8B/BP2CsLzk67+TgHsv0fVmjWAAoHgw8ysGEJwhi5lbqld1I9/ExE+8pLe
Rcxq+CLHkG2vjp+DIOs1ddmtubtc6nr4hzymoSPPrr3uvMm6gMHSvRdMN0D4s8QY
UDiNiOmszMsoppwRVMwuB3m33alv49BiaR/KX5Xo1RsKH6uBydLrCvAD3D7AVrRL
MoLcKhKRq9Y4C3H8SstJ8x9XQ/TAmSdcA+wnNNdfl0yHWHcFVkQwX+dCRCkxvDmX
oUbxvdv+/4L0p2WKdqmmzm2EQ6IscTkn55Hri8XXTzvo7xJPOVqW64fkuWfEf7VJ
aBSmO2IW/qj2u2tf1Mx0ZaSeKAKZQdSxhEG3UwqhNMRnyG0UMiiDTpP26uPgTRP5
JjCC8wKG9fROZmI6E1of94j9V97W9Qpg/zi0KT8x7IQoclTR7yzw/hmwxgX9qmLm
YyvgeFkExmZR92gvcy/pVtkbvq1I7mCWlsOoFryczFexA49GiQRSCFENNgORDQQD
Hzl6xH2mzxRM39y8RgYPm4kRy/Uwvg8zqe7B+giC+OoxZ/A5+nSa5NbFI+Uh/Zjs
e/oqzBtYAG1CY/CQnZNRkYNo/+prPFEvbvWmdkHNtiKVl7uWJkzaoW3m1FO6aWZa
7USGlUd3f7dK74foTwdiCirhHGIWqCfMNmHYXDtHQavjDtArZqMAUmeKcpE8BYqO
gB8oId4JnfDBBCB+J5bb6X5I/IbGfymOgR0uAmf+jRwTYmolhd8Xoq5u6h7g8s26
iIeDkzlT9YNwN+Osb9Ijeb0Wu4oE7N7Se6hWto6Urng9WPd16M+N3g7oUDgantkS
T4yOz5DmWa/m4qhrZI5bMWUjb+l3PafQ3uzSQqnWG0ukNXle4FSJQdTNBlE4XWaK
gLJAPGtMmCcTNEUn4HlvE9gKb0NdjTlVg4AR3INUXIwoakGaw+O9hhWcLipqTDal
QqyznKdHyd/OJ2q94whvMT5Nb6PmLgzfcDm9D/c8Q3EsoYy8rvSaqlVfUcvL6xbw
AwBuXD7KRt1V0+HBxwT5tKkFmd4XOpcPN25vmMJPWmCFpOcbUm43GXbpXF+oapkd
qtq/lKZo5F4XetdHCNXykc4GoKKRA9tQdnYSWkUj+TvES74VCGWsgX4vvKeJ+ecO
KZE+3iqX+wDBpO1anwQGTZLstEnoZ2f/PUHvvA7Gml3BpGlZO01rbIxEgffEzGNS
FmI36ElwAHA4fGI+M8XJDA9XiBobvasW34327STTHi15Ccjhg+UhwmTRYDhxZTFN
LOOweWSNfTvE2Ksuy3Ogb8myAs1aj/nRPKvq+35QiK5+XIo3BpNGrlx5JM+o7nXR
TJpw6qGSkNhavhaUmP3lr2hTfUAywumROij8uhIx+F/QRco44NOmrTNaww1zHXU4
3CytPmdGq69ta1ucCGpOOFuzm9erDvbBZOJm5eaIWi5HT+X0sy3POEY5t2SMIIy7
dMQZ/tzsAwAZSFGW1QFrviq4CKBmsz+TZajMNKnWNXBhIzgP9iiYh/iI2IZrJFQ+
ad9EdNvUIQYBgXzoyIGXt2HaTTsqXnRrmcf8JTGuvgZRWE0Z7su5UrWTnxszxQ+j
frTwDn8Jk1OkNFUnqLVKxUEkP3/5xyxSyMPojun3vZoGfDAnLWWAqFe5zfGf2Qqy
BIpNzrMClgnUjVvTfm0KruwNLLMUTjCOdQTUnS2+DAtxj0/spXncAi/nxLLUKRS5
PQssfOrpfqU42BaDT5OMM5SG/+I0CSs/K/XjJMj+IbE4YXDeRfXdSYAgk7worpf6
Al9fucCzDnAUJPwOXuFgq9KbC8yzYdMJfQZi+7CtwUqMGbxh5tnQ4GcKkbJq8oB1
CRlNX3tXiQS9M0O107CNpNA6MlP2VWixw0otVUiayOpOTzR+7wlGn7EKBgSyvNH/
j3xkpc4PgrqikuZdNTZLHg7Ns9EzRaTLBLCKmYdcrYc9XQGn3Gr9KNDzSeLikzdO
kmSjeEKpvhaObfneC0HI93HXX7IH9JgowX7bIdWAe+AyGj/C391uUWUUzo5huBTZ
dk5ShMB1xC4qmi3o0q9dLKDIuCF1h0bS2XjCZaVDFZPNoQEEWbM+pLZb/YMZuN4U
9VCooq9rEDEYmT6FouDCpdawj3GObkaJrB8bWbrGnOaYIE7YvzrfoVAhjervGgeQ
skfYP83Ow5u8cIVZbynjP5rbOxEPGfAiNUOt0ROPwieQKy6+e4VR/VSuO/HGGhfv
v8Y+g4tqrcKXsQ1ar7acScj8eOSTZGGRtsWegRQYFA19ZsAQHFlGDoY3rw4FLjOy
T6kYrbELS5h97zz19ztcvlhz8kjvZisDOpiDiiFrkk1WdcJyxSYsCR16RRKP8trL
3Jl2W+vNGs1ef+073rbRr4JUqr08cIYz+nZCpoGO94Qz3uh3peVpOzJQvPqjjHq5
rVfitT7WOCbz9umnJJKwU4kucgxpoxXbXq/2L8pNSnplAHY0LpzsiEdlXyYllJip
IINeaVmY25wBFdbY0VVIKTCZwUyU1UMKPGZqv4fZ0t5odGYx3gzTLjnCKei2ca6N
wlikifvL6Ksu6NJq/WEX+a7Kcqylmu4hCFBAwK0m74a++L9ubxNZR0qMmxLvInfN
h7FxoP9HeYYC1BDd2x/7qXPba81L7X/BSC6N7j2FQFHJudZo+FZv2i5j2/mRTewI
mPtizWMYuSaTAXsJ4Cn3uV7IurRtPAJ1ssd5zi8kKvoU0mlIZe7wwcsNDyxrNLg1
M+fIxgBze1T3y6q0Y3rF1Zp48WArcQnuMA3VV10yYfaUODb1Ve+awFmrxvPcTucB
Qarjtdd2pwXSL65Rd/at5PQyTAEZbTewLlnv+Kb430szr0sNyBB8D+yjLgNQMnv1
CK6p8cLBTNSqHIssF6I3XXMiM/sMr9Ij9p0dQig4cnJONZgpY4O2ZXMXQjK5JeSb
q0W5yw/5DQU1OH3qsDW1HoEB9++NiUYx7GfejnjldBDfWdU5qnJJ0rh7TZJvwYH7
U1VVQ3aE7piqPalIpbL2wY0IcK/hA6wsZ7mIIA5UghI23qg2PT+PrNbvvJt1jF4g
Zg58ip+Yr1EOmcAyz28niMBvw6E1Uki9AYjFD1kXUrm34km6etWsFVaFC8NEvBBx
RDvXJzW3w1E1dtDu4hem8eYmDPkWmQTeo12VuwqrYEw0pCC99A0Y7JVEnm4XmL0J
qKqMmUROfNg2KfZZxJ8p5M9vapTaF8jT+XSEBBlIcKN9HmcelcX8bM31dhdeyFjr
eGqsZzTIUlEmBnghQj/t1SBDQ0VCubseO+UyfPnwaQULofCD4Oq3fIsMQZ2UosZg
b/rhU5r+JAobTw5znWFx8lS0cNg8J25AhwniwW3Qi2Pbl7y4lMtND211bOsfLo9+
xeyoXdINNHVEK8J/nJKukhVbgHgkQ+SdMe2EyMY1gd6mkaBkKc2FY5mYMHPJbzeq
m3PkkoCxGAFHNc7/z6hiQe3D/5Qq/4Q3GTwMtt3nduzhUOrcUYBvF0H5lfBCyS19
imp/jd++bmX/nq6XdDvW/2PKV6WPtJYRhRE7j2hQCnoS/CjoTH9DoJ8KRP7cwiib
8uIb3bXcMG+ZP7sIdBg6GDR9n1QEJOIQeBV1ifiSJgqI5Bd/Dl02DJbZq7WUe1VN
0e5y7TmtEfm+NrPpC9Y0cHUGxEvzO09RJCt0+jOEmkGkw8iDaXK9ldOG3B5GnR6P
93NgzcxK+RDaZCZ2V6oqNth+AFvmTC4MvWXMoUCmh0A3IwYrO6JxAIB6uNnQYhvf
bAX00ZpLzfnwyJPa3NWZfTZamRVDVdHLB6Rj02V7uLHqobysluIGPrOEeKefoZoG
klvejdgjkzCGWob6bqiXqXUewmmCiGcXF8wLM4FzMVeO4zVwm/jXwVN6nJDIWwcX
22Zgi32BBhWGrqHjcaxLxoD0zoj6uU/OwUtQAgqdFxIohUw/VovGGSX6tw1iEZLd
3tCcfCfIQKfCxLGAPtE4DAsXuP73O5NNnx+uUykNGHtJ87FeAYVirzonO4ma6WzD
I8PlCRB+nBGKD+LYtE+VMSTpZz7wDPm8dCIWCQJGpLSc5jQCD0QXK8n3hkvGgLIq
rjTgDkjcpPc9ax6jeOis5Zw85tXPEiJpe4SZQmqVR7z30UvAz5GQhNSoOqocHUgh
P6lRq/1HTBFFz9ye7R02ucTWEnuigNFR9d7O8uQYxVXXYXIrQ80FOVimDv4acy27
n9sb9SsU9DQYUwuWRisfFDxcWKp2+PRYuFanzdIQIbEhz/a3B12yQOjR7RSRP9q4
axUiLcqggEh+WxTyhGt6OUJXw2U59sSmkr/KsJC8n9xTwGUnHZWVbEehQv9H6Uhk
5cZAriYcfyifbxUV0AlfiuX/Ip4XZqp7kU/BH4MMook4RNYxgbLUJLwV0HT0d6zH
9+z2jOln3klCl3ERPL6vC+4Iu7mgvy3P7Bas0Go8DghfqQl5dAo0yssb8voWH+8Y
EUfdAwHvfn4REpF2LriMfD8gSx8hMKDOnMIQs+qeU0IjzJUTdJzJZnHiLMYC224D
SBs6QQulT8ven0L+ptLltOaWdb3Sp4ixaGSvCTtgrZJzFYaUXbnIoAi82vRGK5fP
oYzVR1kV0tVKQarTrGac9s1NoG3qfoiTXkMj+5pJvU0rEtufLtq9owkENsowyuJU
6J1pB0E+HPquTJ9hVT9dlfTL35xrMwTxiiNeCNCNA3Kt2rE3g8RFHM16trJIqEGG
ewisgxDoD/M6VqIQcpesibUj4vXTHQrJ4p7kK/dmkhD6hvNPFYl6E1585sgjCKZA
6/HjoJqjJ/ReZetJTLTVeXkL0y0vnKUdHXRhNQmkEdmfQK6d3kbCcG/Bh6f/c65D
UtdW9jIUrl7x9HjRMhfpFsevK4N3sZR4dT2A1s/HF8VRpT0JsiW53hT8ogC72k41
Q+7KsKdHKVCAeRPam2xguQNd4bzOHk5T9I16sCJNyCHSmZqgJqCjcHy23R9r2C5n
Q8sCHI/AVBymvhgeKGWZ46VOqBJcf4jjkuU3HjmQrhOiKKE9qVesVulRoBzEnjWo
7LNSHw56m2e2bI0Kp16qJ8b9eA7PQxuTgFDIk5c3FPSGZg3CNrHkOrOVh3LnMMi1
jf8NfTEYWLtbMrvNm5C+ysE1wSncJ27WTvzQtmHT6D2ndeOrGwtJTmj5o0GX0f1K
Trh1anlPVyLqLjajDaYkqaDxqP/oJULBLCGgZimJFF7Xipy0s0l50U2b35z7ZJK1
pmZarG17KcuqFg4vYxU2p7FIVl307WNuTB6AYroJwVXLyt7CVhXSrwcErzcG5tbk
qXoycObkNIXlpu4grSZOkKRu+2pemc+qAJpNfgHHbsShSai0Eh1L83fm86MVUZg8
tTCb/kycIEFfzSvobqJt6x4rYCBdvxpggIrHY8aMTIIV+3W68Ueps9oJAOF4O7vZ
eGZBd+A3Wp8+VYq2tk6PtVWkIOdaW10P/2MhRC2Sm1R+VwKOg6BgZsTaCCjkGJqy
DmYqgl2jnO3ErtjfbeSQVB+nyKI6142zY0nEICMOS39ytAvfQAJQaqOPhUCzhrnE
sZCtiImUQs+ZEhWlIHOMu0KoYsSBhBSKBhljGij2JLg8yAVijvT8QWGYczpwP1Fe
gPtTSrFbTesxddhwJiD4wOpyRHirDEC9tLLfL5hzrJKsEKA87yWSHDzTNT3+F1aj
bRp25FcomIwYYhAImC9DPhukI4yJovmp+U5+GgbyIhIXQBXEfXGQJ45NI9MVWYrZ
sTtFp0wNzERKBT6swehDb4M+O9/phWf5AH9hPjrVc+rwNT2gDALfcbZqerXrerfX
c1VmYVwdo70pylDWRr5LWNZzOwALCw3v5+ZcuoULRNJcsT16tAC2gQT+9wToH8LK
/7u+VmBBXi6aT0S83SGIvsp4P1oAhyvnqkuoUsCk8StMwubBvGUELn3vqingYnaq
PgkOxWY7EaTOa5W3JB7c5N2aovcuvQ1klQL4aW4t3P1dohsMyOJaUbvK3GKGqN5h
wd27L1vE1cz9cx0ARGoiM9YqfwGJ9k9dT2vUUHWi1bhpGROC3A86CKU0JI3Jmbku
qPAs/lBFEq5ixzftb0UGW7Xh1vD59nPRsYucmlQLPa/ZRkkhH8CqS5FRGWHk2BT8
Q/y6C3hEpe2WbTD1rgnRUd2pkIAybc2O3GDpSiZAScTeIXrjAEGYGahnjpN7Rarx
4+IwRrCcHddWxtr/iJPJryeFo2dkPGd5ypuefGGHhu47bTTbaF94NLRk5XewT4f6
XGLoixvf5vMS1CeVRvDOYFPQdqxNHX0kpCjIo2+OPfHbusmRiUU5faDv2fZTu4WO
vgcTIygv/fyc6IkSgi8Rq7TOV5Id7LEVhJdft4vnAnWmQlRKTFYE+d6hIxZ5HsVS
8IqEzdmSe5CyDSDpxo0//U9HMytahJcdV5AbYpE/XSCS5rH1jy+Kkf2xG04mTOKB
S/iZqXsYt1o0BGhGbVCvLLh4dAXGokEa2yWDM4d+Zr/frcT7+RdOqibbT0+7QG17
41PEOZeOP8NGahE3ScIfNqm0tGymCq+aJm9Wt0NDA5YKnSKaOd4hMhHiovHmeZQY
fR6nb+6aPQjSzmvrqouKqN72lmNwor33tS59ayAISjSQARuUE6V9SuSzOmU9+rnR
AtvvsS73QCzys5SqAwWgH9NXCCaLpPP513oJLwD4fWOa7BEwjhemY5X2UuJEQHng
8AOVttMR05hGIvzp9wLuQRqZEtTDuwlGZlrG47SUJfA3mWerVJ4iPOSjdDMNMMZp
8aIiCUzqorI3OPjVtrxgp3c940QicnZADHktHVE29+0qS7R0BPHzHCqLxX746nND
fKbQ2HjV82jFZb9RGYZMBjrPbveeXuvOVUmm51Lygs+LidpTPLIcoMrzbzgb08gu
aaeCQAMaDE4RVhzyeLDA5BwjnbWJLSaVqAx1WC8o6xF0VNUNiLHH3upPccAu5Ud2
rhBhy18Z7WLcjWJFWjg2JRALovvcTN5awuGgj3CEHkf00Xcz+plkOo/ddXzp2GMn
4w/DcjwZbpOu+c2jsb/4KlLUdi1NbqmhejMpY8OjLjUhZ83Pp/k4rKESo7/NdJd6
UqboEJ6uaG52r2WutWzCgLA7NeaLGsk/2/WYy95FFL271UPKuxb4pEXI5zrZFlgU
5VXgVgzrIsKPa0YvIeKYA++dIa/0OEJ+EekBAiPJLVeOP3hidhVOIv5dBDuJ/IzZ
rBnLgs32Efe+2QxxoowKnjj2f94svp6923sYDlc8zBCii6yAb9xhl1YtlhzjqPBe
iyxRtO4OKqoVlAl0rK8fnaITZKTj17tKCPGfMJBcgcsPFlkLY7DPZVa7CJgc2tVg
7JA7gLiY+j5LW/8WwEvY6qsY0fcF2Z00+JdPPT8DG4Rk59FFvFRN8AgpABerYtP4
EmmiLz3/Q3R2ElJtN/9aIa6FEqhSyePQRT8+lQ2ne5TkBWwqYOMbA4w0KlGuPN3o
W0ab3uZuAJL+nxTaX+Bc7iptLHLwmQQ06GGIf0GaDr7ad5yXQ8KuZ5xilZt0brD0
s0MNariy5eNcxIjAx5JhuJC5ZGeyBF2LvF21deao0KPi6nI5RC44pgnfWprrl0dQ
uY4084GOEHGPEE/jkGsMW+DM/O6y8H04SdZAxuWtDI878fXpJS4cJqiJtGSYfbPy
9o8UWVLA1ZESzKxx8YJTvg+MBMKwopD94+8+iuYItVVC1JG8Mynr2QWso2eyxciZ
EBBXrrIzrl/gH11VFi6N2c4QJUcwHbElaTQHfkYzF0Jl4PNZVigU1v5hE6aOkGNK
HsFEWWrQ3KK6wDjsROn51LuLNdo78gZzSxncG8TuZD70DKxi2QMCI1C4lF7UuqwY
CVatQOXQPsGU+1mwsXubrIamK2KPihFSyvCNx1OTvfSXc8l7ENOq5X4ZxyZhRIAH
gUYgO8PJNlh06SEZZcT9FAlbmOYnXofvhJ2Y8L9MU1ERfoodm5N5yr5fBu4tV5F4
BS2BlxrQr6kS/XEJi8cmpaGcqHntOaByneNoCjb2sDHHW2ShygGTXOmSr4N9i3pa
iCP04tuiqjr47VKLOvd279Up7kmHTQCAFO6xBGiimTwOQFirGCH3BrNPYXDNWJk/
i18XO6b0dyDmYrHjABTtzyqN4SEfbZjugNP8KFTNsJGDtn6h1G6ljK5bu8Xn6MoF
Ows9hAJYalWSRMRK4rIQ38TssVuIyvVFBmKiSI7DB7yB2+rbEl5fXFu2SHPRN4qP
AOIM7ol+nTMnBXdLssiSMe8cEknu/s2P1PG6ZVF1lJWv2SwsneU6UirOO6x5NL+/
GpnPMseS2G3Dx9Id0JpcwG1z3BC6pXZtg2AqFgC68myNheU3dQr713Xm9E4PVWom
f1abVhXth30ltbs7O4KKP63piUA/RKBigGwTlBYYRpokHtr6gcMQBnq+UnxgaTFu
N/Ruryxr9Oi7KdcUgPxz1++gO7+O4UHlZ5G+NjO/qaxwVmluXIUf37Gv8BCBxWvB
+TUzJSRTLuXAT3DzFX8TsMeD4Q9wM3OJ5PAjJ2YgfeIA06ScK+PDNoON+6lWa7lY
2ulyJskfPOhS3wvXeqweaXoQAOhHWmBrQDVjW9dZ51lRfxhxHbyzySeWzZPv7GZ+
POTW2Z65+T1vptDshI8idzcaE6jvM59PQxOoRJxzjxucvuZ5Aw4JsiS/L+vCHmxY
Ey2qw5a5Hz9uKSX3y/7sRzXfdxh62S9AzH5qYMYA3RbCIdaSeQmQrZ6hysLsBcCp
DfMhUGw1VPoimK4ikWVGk2dDHhr5NsbaWTUxPLMU2gLhiBDC578HUbCl91uw/HWu
3JIfwAdHhTMuuM8xuNHypzl5TzsBRAu9ERv3ZB75uF7YatuJLwYK9a0mcR7tliXI
AIQDlaTDA+o92oH5DB682TFh16eFF7EKdCfk+j4mI1CmlaQ8eC2W/INQg+l6AznI
cZv6/NWYud6LUfJH8lF/OedKUDqn/XnLLZy8p2MzW/jpGJWQtOHEO3RiBLWxtuBH
ubLBt7f+6yPhK5IDkALWV8/aMTrva5VeQOngd+D0jvGWdi1+MYjy90UyBOh7ewJY
rNhbjd9oTQ3d06jS8wtZ9tju7ujYdyDugNcMe2j3NV5Bllf8ZEDqGN/q4nijJhZJ
7YS2COgp7FzOuS0wgcB55xKyBUeuQA5WFjYVSew+5zV5xjEdkfHtBt6yA6PgXD1p
VAVvPsNOtSaFGEJOrjr7FgL0Hp4SD0n8AtYPQhfuRf0QT6dK0oXfqmxc7l9CrCBo
D0mOQKGtYhk7IwIpiyutlEZkjQiEKlBGZjfsr4dUgNd+OAdtz3h+O9OUGj0qV52n
ZxxGE9IdokdEBW0Yg//RNG2gjj1IN23sW1A3cTqfxbArZhscSXxM0Ge2zaiSZolr
mVRym3BtMbsfIpndUvslCqJooK3r/C0QbOjPQnpfmUH06MV4LBgV05c8CUTXBJkr
KEgL2n/ercYR6hYi9UVFJ7T9gGnTshlvvfGxUVcZQd2FlXlwEc+8aa7OchD0n/Vp
WU/FWuIJ5a5s3DLw00L+848idAXLbQgElDkSMwy6GervNS6sAsL7zVgClO7b8r5C
TVSfWZwZEZzjcd1dlcoa04Ei66uhd43ThYBUigmgypil3oM5xVqDTzXkQLtj70B6
Fp8e0nRlcFEDcCh0eH4/qBpv556rZpqQApkpnLUoyWy/qRBynkx/o0hzEXgEYyqV
mcdWRVPwWEOHLQmWrSfOXU6IXBMI3PC6z31XB01yXmLSijzxIKOQJLZyuOkb9qAk
BcCjaSVfaS9/gfgHQvQZuzw0xAsQbxKtzby6lsEW757UeSSbDkqtL4WbHXPFH61P
I4tivTt4GkON7cGDknO4gmEOuRdNg7Md0OhwSpDcUsQWB09dYF2ZGtoavTKIHpn+
ktDU+YYqVGB4rtZeKEKNfC4Voh2NCywb7bdp3tZSNmjzsZmlzyelNCJ3Uxq5q4oQ
GOhb8/eF1/0DGa7VLvl0Y1ToP21LJNR3v6VsDyMfJns9go012KtTEJGc7J8QQgaN
Dqp7ZGM/+/4e0vc8XqHM6IdKzkvymveni4JJr5EWOFB7P6IHLulFH0ZpCIIVpG0n
9je7/cLR7DeoQI9pNEXVvDuZSViNJJFK8OtmbnAMkkVzKqVk4EL+Kd+BLjjaOoc2
NRqNsr7OcvKg88VPt//Fi5tdHSJ3bdEddmchH3DblGhCXdhbQw3I8ug3qZ3EqCbs
mFl8ggq6w6q2P8fibPtdKKl/TKM6fXcMja1xXMLxkTF/c70/txqpRHEp7KDL/rQ5
iJ5owMRMAg2SULNM/qPriSstvOT5Z89ZnYDiMM9jc30fpdvynFjbHbjcgmlrrkZb
Rfyhlqxw/acFeObvj+gbQRKW+PcEfao8vS3MVXXsTV/bnfxoW+jBOIzrcm72OUtn
9x0gU9OIl6GA9UdeGKP1mXolH8nYDrBbN3DcubnhKuowx5c1rATAnniXoTE53h3q
4PzKp2VX/5PB/td27NzDtaf6ig53mrXFT6o051YcLel9ZDiRi1Utt+uZcVgtry+p
PCN5awoyyA+x/ZjixcOztkSl2EmvKNwOG3PP496WOhlWzFL6B6lcPNxwmc8OswbP
9hYPV1EE9Qr7BTMtSdiCMrdyw0F9wejJba4be/EyVVeDuDEYX+aL8pCDuzX6s3sG
078MyhdmBhQqoWIZrbdapGw1gh5Lr2UG+RkmqBkEOBzKdjsp43Au+5y1wGCWv1Pw
IUF2s5NP1BBuqqW4nGgMpSptsLmVZIv4NZH6qENe/sGjPtmhr7lHQDGblKGloPW/
ff7xB8ovLH28SOerqpOMbwGs4xdCsESfdTFpsDnysSNIsTMbE0qT8QdutXZb3uAF
y76zLJciU/gZKilsvjTmih0IQMDLbKRfIGl8ylFmfwAt82P80S2e4wXrxDono/8C
EpzB/e55DQBdpbT+mV+6++hfnCRq6R9KOC7mhB4gvW89DyouYS9y7BrHNhZR4OwV
FuaRTPdXjJKsn41YAhA18s7uWERZsALs/Tt6IS2T1DSjXqVpEY1EJjDB7GIBza3E
swAPe9oT6jmis9xyeZVeiXgc27ZbhaTACoPSKFcXq3hQ0pZL4X4sNdKlRL4aqJur
hDv9yk/AGZNfyR9MYzqQ9rFGLeqP0kOD4p2fzg5jQH0MBId6QVuxLLylShxzvG4d
gRhXyTb42DagAeQWGAP0MeHMMGjncOTt8u+mkgN7s5+3ei1UO2czJuIhoVb+6Dcq
Ua4CeBplbiMOQqHBwhLhHy3vJm0XNhN7Bcs0YYkyaLuxnBRc6e4pewI7jCf5Qcrv
WJLMcI+Fm1znNGjGwkEmBkS39bnpn+LJDOz1cjwIiEUD5WyUYfFIp2/X3G35jqtd
LZp4jSi3hXCK5tQgKth9NE3wyy6JlLdotpjwg92NPt5tQYZtZR2DVP+BRvuda2Iw
ULYLHi5DxFhjrqcN8cVmX+CwFsScTBPGGjONp4aO14XxKgQ56u0qAK5Xiks9RUXz
GVDnSSIz4K6s0G5kr+CD50mRgrQXm2DoB7hOdNDNWyxeUTnBUSLnfpTYhJ9j1OOJ
u1j5s2wbaRJho39WWkYXHioZiEyJGpTH8a+J/ql+H+ma+ByCEsXPpyxuRDFzmHvH
8X9cU2MtsuvqL9jyucjCLt19s/K2dnV9zXNX5BOICjMkup5R7G4TaydgbHd0KwAE
7vEmcWmamfHtwdMkMZj5NhAonCRQRKgrpteO5oA63vEPJr2fTuKnPpxnX0ckgMAx
2ro/DA/Q5BGMGWARaAwFvW04UeuKO9NRPOzG6xrlC0quUwPCAQfeveRWtQW34s3/
L3r0YVDyNCu6QExNxlCFdyibisMOIWVuZs4ssnEDL679VsWvSWkd5/amuqm2FH+C
Qme5wxqPQEnx9vAcvpj0YpLRFwV0AvBWzj1VoUW6Co6X1Jh6pSdyUusB6htrEsW3
HkSeHsRcU1loM3QwyUq7rpO6AkZiFJ9oXSJH2HGcudChVFWW6omyPnHSb56AYTJu
ysnd7aDGW9C66EGWNCH7WdrsbShb9S+sC9+dRs4/xpXmvBfACNlPU45Nep4LnXk8
xB7q4n1wp5P51uwQtZDy8TwL9ksc9Z1UlBcVcWs7NorRNnE5+A6Ei82f1S7iQDrC
0OrJ3f/yZNh+qBY7wLcdPUm86HpntFLGJNmsjqQ2AgxguV/98xE6PDx0j8cg9Kn+
F61L2MYIVAo1AUBQe6pIMxV0BZj8aQLez/MlL7uk0u+YQapgEc7jiZyIadOhx6Cy
MHCZWBoCHKzc0MhawnUhXG8G54M3xAHvdjdoBBbH0/dPqvtgQHQXJDD+wRRuAoB5
vSGhJBfgTJyJxu5/EjMFvt95xgZy35F4dYT41m5Psz85TUwZGzYlJYIePUxonRmk
CDZQDfqjpfnZErk4YybNVJ+pHar4RUmC0CMbgTbabTIKL3DdTDIEXCUUv7qedrsE
dzBchagE0hB6/KQQVsGVZPeVQHOw0v4EY3hsP7eLDg6nstULbSkhCw1sLwPa6PMr
Pd/0Hli5h5oOQc22ozgg60nb1WNsFVtuszi8NWuVD6Ee2Cp6ifQQ0iMUqPHK8xih
Djs3iB9OX8LBVET6HXP4pmogHGNVNkI0sPo1kJyXmmTN2B5tSJy/7e8ViF6VDQXS
6LSd0vEaOqO9iB/qP5mWTp1fu7l572auLCAZZO4jweMEfnEm3/20ncQv7RMtMO/d
rtZVubRdP4eE2iTinBwVqu7PTOyXqUqxlooi7yFxbZEf6nEicP51bYxYIV2Bz8jH
3pqaOCY10ZyAStdLSpUlDGhI5v9civmpxqDdndHAZNcCu/W/pNqKvk6DtzaJ/TTt
gRWeWfmqhBwvegPm8VecV9zc1CX0i5M4YzWhSbfqJe5pena6HMSLcv1+tTRTCtVi
aNBca3kn2+A1dT9U1Qlqz+9WWHZCnLnEJTzv52R9GCrNFkP2WxTi/gRxX5gg3lQM
Ds6cA6mm1wahvMgz11BriFXNPbY4psf0MgRQwFXYANhQKtTqxQJmYCw/AvbHhUCw
CCPDH3lVV1zQXDOD7SnznjW60SZtNAT0wQSCfaYohzO/ZkiCop6wETFZHxmUO4Go
IpYkVtLaA0lSUG0wYhQSGz/YSZzNjp7YEDvYnraZr/MaJyjAMDLS323SRIkqnfzp
fTQdNflm5sJDeYNKwLnE5SThFHr1ZTx6CeQuEzn6AloZvdWnnXd+fGwd/Qjsbhlt
uu66wruPDPC884fFS0go9L4kyGMqvGv3Q+yP3sCuIYscPeobGlcIZoJXKzBpV4X9
jdFAqGtsTbnbfDROifFBETN7CmR0s/RAtwKbm7FBE+dC0FVWlGiVhQpMQWcI6R5p
OgD8WOc2+XunRK/s2xkKFu2Acf0H/GvRh20k49TliPBGLCLZBX7265aSMN9lZwkL
MqNVrvs4Dya/86aIv0EDh/hntG3ZTWx8RLUnl8F4AZFziCURUQoI84T2EpERw8Ma
Xp07bPFqFMaGbtJAfqvC9IWB9Skfh0EqHyKj6QUMieRoYwZjRhbo1prdLN8Z5WzM
xWQiS+5gW0Ettld9ltNrqh9mYCN/TKTgMulQRXr5wI2nEjUX0/mRXM3AB0u+UDvt
EcO0RKepy9xmeO2DLk1INzVOx+6z1OAUiaC5u/DV1rPqJfFSrA9UjdAn/UnkGVjq
i6P9PfILDs1Zho9qV3fvh6mgFyi+wDP2yuvw3d5nRN/cEICmtVx0RvHd+c6jCRx8
V5S77ixQGo2bEaEdWl5fXXacikXYu0fpYHnB8iUiDqFdWUVrUOZ2B/1WrtA+wwvn
W4SUPaTNY2L3yTTg4J3n9MgVLDXVQkuRwlFPc/Xb+aJxVuP03HErX4WaBV6QKlwT
v9aNESZhgeoSh6TCZI+Esle7QpKA35IoctVtbSxSmudRZ+YJ7aAZSqTNGs5pOIyJ
SAzeJbs8LHNFACwLkrvqXECT/pW2BntYcFq/QwUiowniRvLlpo+mdZWnF9IeUpRA
hcvkDf7f7gd6Ws5rhTGz4hBDDhBRyxX7cymuhZu+uc4OC1956pr3xAWEZvDZKqED
dhLA0IvTRssAdXcwX+GRInAwwM2pGjiLCvP2ScuIZ7Tvxi2FR3nR3+Q15kAwshBP
zhVcgn64dplf9ab9Bflc7h7pRQAFP70r1CsOJu0CVtG0f9C30ppXSMuE0rSaBRiM
fHxXbVnnQoI7dXj0eZxmdlSTxr2mkyKZUoU0nJi14D8OhP3HG/oN/4nlLcHG0B8D
W9K2Zyjp7jAtsC9Q9zpe2/ugtAN1JIQ3COEv0CUkrKHB+hM2PbU1AeCpoAoU6INp
5u2+qewXCEpqj+kBwbVcIJoABhy806Qkr5r7eR22GTrcYgNmqTPZXZ+U6CQ6A3/q
3TN2RKdLgOMP6VOGkoqwF7rXqGkHNJRSLLIFp+c/fQP3eomOAaBppMD07YITnUgX
uu+E7jyHZpysH2lfT2JEjOVnUoZ4EVvzTsvek5o/C0kNQzoy9v4unELGykv+yKHy
yv5o6ld1PsQdgClRJlahQSOH0DmBZ8mdebQzMqcsILhxQk71Bw9Tg9Cu2SIZKp8k
e0braciogudovVuQawfHaHbqy7/auLmJ0Cc1UvGUgu2f7MjMhvneETlUr1HJ12St
ckMKkyS8faVMn1QtF7mXho/VRSeVJpyXzDq7bJSp12v17uZ8HF+Ft+dhGkdIXIf2
S4Pk0l872M1DPdXY/pwaTTB3/fiPapgACQPZ6Y18+Qe/xF2YXEGEdyMD2sfLtaT1
y3/xXm4p4Wlj8SAMd+KnlbQnTqGm5VJr3grTLOs0oRJbMZyBvu9oPgglxUlYgRq1
vM3ueqbdL77RW7GPba/BysRr+E3r25EmmPZZgGMj5lFaKV+9keMzHvCi9j23UjW0
1HFiCQw58sZZ6IF41Sf3Zne72UD9tMyqzC4SPZHiX2GOtGTnzjNFNhUB+bIAlrAm
Pt+yvyv7QcWhSseqewKqrM476GK11EMAU9gVc7OfK8ETbOfc7FXWEVX76baOHgda
f49i/VVwUAHHql81WxIcEL/spVHG8WGuRt10Hulp4yjnsFfSDif6uCnuqLXneQms
XMK178sHgsv5S0W9LP1V4188nZNIsIdAwNYliuoV8AMXI6q/rJWeKrWRys0z45hL
I3b0aujHiNq/HVaI5w+2qiwsmJ/777zm/jgXjAoN8gt1SAV4979e8sI/DJFJOv3p
3ZCWiVje3ydeeiP2RsAGybH8w37zxdY6KZZ1qyUUG64Itsm5XSSCnBpzArqYzkyg
rrHsSaIDH9RH3uZCq33hyK6X17ItzMrWlNg5nSRfZT5b+cYfUvS2Ca2Ge8OfZXtF
J1LS7fQwAmmGM+kokQZtDndj3EkUU2mYBITXyrJTojKjsvEWmtcrsAi4sAP9v0MG
S83wzE9aIu4Jjj3RDmkpeIQOAQ9NiFleTXq5ysahfdtsr32mUPIJgTNLAu7ibCl2
jiv9RuA1BtcKWeoJtFee6r1kR26wwXaAT12l132tDPg8RKFw/d8LsMuusS4r1Zxo
K3MXYkurT7nEHGibj1vQkZwglLXFxeSMoj2s/IcyMc9hzDP6C+kS3KcqgG9uEKLC
oqbklsvCHIi2qa9oTWHx01ziJ1vQmfjBAJcRI78uaGmBqvc5ACi+ivAYoRyvLHJ/
fqgB7NpfbY1ZXrwuWZrcjv0GV4Kgwctx3aHk1nxJEA1BszmkSGcQqu4aqEje7eYb
VZfaKSlGe+myJ7T8VrrVrmf4qv1lJpoUC3L9DiZxbVLcPM5GaCBk+NjT1wQyew3C
DIvvrpnwZtcevOxk3/JkdnDHvDeLMx2YjrKok/Ng7BKygMQzx6AxW2T0rqbiSPaH
u90S6/ehpUA8nhrB7W9MEud6dQtOk1yu+TUYDrLSgLZW5ebJ19Cdcxf4Ac8x7A9I
7XMi9KmVNVkTkbIu/qhAcwJZMO7BEC97ZgoEL7Q7BTVISxcZXgv6aB9BBNw8FT+O
tmxU/wCTez97SKLsJpBQf3BvDS5w8a7VZWoRGezax9OnFqXQ9g4edtJr4cCWY767
JaIGxz8nYI1VZd263AuoAwmA22v9N3Zhv2BQaw0ILredgtitv547n3lJLm6puvC+
NrSqvbxKmycJG2sREjfXksz5LKVZLQ+cBj7Rj05ogB2/W1kQczg1WUf9yz4zQby4
K6V62QFp0HLL+6d2N7w2D/vk2UJHmoVMzZKq5sCuE+p2r43fsLb5OrXH7RGYaQb2
+CzSVF5xjjByt4w6dXGHK2K9mw1KLZhGsSrIo4oBX9N3RIjy9kE3MDx2A/HZc/V2
CLYsOtlpJijvQtGWiYOaXU+iZX32gHwi8h2oI+0UCECvTfB0Klb77I0nqnlKoIU+
me23B8QRwirbZJgJiYb5dSWymr2Bxtz5g8aTETMwtoTuViR7irEXU4TSEin8BOCW
0k9ZgdvO0KdB8JBGU9v2eOycSpssPXIontxRZA6+OkyoxVAhEmuOgwEJbSa/d/yo
wDcHPIsVwgDOZBAuIywUVlNPPBIewQas1HL4bv12JwuHCdJYTWBaSTRClUPxFwbZ
jEbrQDkBHr2qmsfeNgOZsE1P4pgbVL1YlQm7euAw/e0YAZTxg03J8uqmaK2VJ2xb
cGRz8syZfwyj92RtYImFU6RJbrSgXXxZ9KJlJgvfYx/X+gtPgD8Cc9SblDFzZfIw
JKkXeR0shBsGkzJqN8t1SvgYTxiEAIdp1EX8Bhh3Oy7+iA2OB8SGGVM+XBgCYKQF
PRkokiCWZNlTE2muRH9xycveSWZqycQ3zwjSQYOjRYco/f0qgdj7ZpV0WxIRH3oN
ppiViuYNhAGiCEPRw8lEy27M1fCwDfGzrhZO+Cqht/QGvD02Qfp7SvKKVH4wxDsn
xAccaSoywyjxBcPCjDErfSgh0bG3fTeOxszFoiYErOpjI4Oql+Pg/Ehk4EGUJtsT
QONseY3kDX2DZr6JAaNJbVwIitg8xmmJh6cOkW1CFm0Xq+qYDIFWw/V4YWUSi4f7
gEUtVQq717NjMlwXnH5JNyW15fkPlmBtJNAbJ7HYNjqJqx0VvpQpc0K2iiJ+KmZC
g8zw/eUqX0n1TudAoWJZXLJZ0PSMNdnkCWJvTbK7diW+dop8UU3ijCGj3ViCA+Hz
ZvDJSE6b5Ejj1FpkWS9oNlJ4pxZpBbrbvgFsUWBnjzHkUsZ/YuoNOWZzIq4I8lph
EtG/dchtCQ654Xx/8gf7NLo4Fe7Xq9Ftjd9ZRVFA9zV2N6GRzNNcPojtSlVseM/j
9RsaJs5prOedRwT3xZ3u/pvgsInMjpNdHx7gzb3hpw3b4PdRhDfZFsuufGJ64p54
l4Q9dIJJklP7DpOvm9RN0rdKmdcQyKr8c81yFStpJrQ95KzA9aIKB8aWplzrsQax
cKdCJm7BKYkfn/ee6tIx/vpgJJWbfliPacq0P2z+RnPdpVxw0dAFurQGBn+iz1sv
V5ApwbiCsar26QkcKJdeTdzXrPkhQSfflzLZl0Hv2D07l5qQXPMyV8d3bHYMsbpC
Qb+9ooGD8VouZQQ+N4JkCJH1AvDxR5OHv/FfR6ZY20jlKKk6sJmji2NBFZZ4Jfx6
Y1ECiJH14wA1PlQf5EE+7AZ2hgEsnFGMp/AGsSZgA1U2o7sHnfbKT4uja8XQghGA
uFsdsJmPUG73nZwkkjHjX0HHFR7OBDHkarhEqo7jNX1ahMTG6xfr1hidGHNTmDBw
u9hswdpVYB1Gun3LO9oXLrJfZ4nlKOAEqJP2FCIScLe13CZpHdaFCrYpT1mtj31Z
3SRPd6juWHfZYxJVgRyLBw6gsiZnPrF5lXShp1M9UEg6XEWW1VDV7YPdqwn2bMr3
FZtslKWWlRp1V/qpUz8VwVoWm/6sIrCz2f2releZB6lz/HltbYgqAJopnq3CeFgV
BTDGGNIIY2UyqA1LfILrE+tBG31Yr9acyY/8AokyoYdyA2uNQsABLZh0Y0fpuNG0
s423mw99wpc3aXI0mBXHC5wYDPj1ElNE3bzk0TPTL7W3dulZt/nAbrH0O8D7B+LA
4Ury8wxXycxf8uMWVJqHcObPWt8+J1uaZeBGfTy5jsn0Wpe9gH1iMwRk2JJaSZp2
ZXBpeqGRSJSQfnbcwsk8kfGvXO0HmMDG26/mxP4BYMDayty+IUrlkI4UHDwqrqOU
F/TXKWnGWTIXsbziGY5124QgvZNHR2ZxBAgouo1Ho2mbQcOtN34EKM4U/V5Yncgs
TT1lXDKTzfwWnZpTcIeHkSaJQu4MPlk+JvCZzDFo5xtWFeP72W/qAjs6+dDxBqoB
2Iu2Ud9yGo5BXseuDd+FjGbsWsYlw9REoXt3Q9y4FlRavLvXmBGSdWME4Bx7IVN6
uMVmTuY0Xp/8kW52sW3lxt7dAvZgzYR0GpopfoqmQ+ufTZUVlTPTtbndgZtv56q4
0COJszeZfS26cVHYgYUxc4K2OBOklyzytp1DZJrr03wMYdYV15vp00arU03J2eKo
RmP1uh3l5iYziqGzU5OwgloGvDHl7puGRMvuK3emWFjqlz0lvuGQmg6ne7xFKZxW
x1sKjL1e9T8OFdhf8YLcLNvMU4yhbVeX3pGFqzIIB7Iq3kSZNewTq/pH55tlAch9
OfRwW64IOJppUtwAN80woABTA7hVthnpMwksIc2XQA1r7AzHUkdbClfq9pdBEhWs
AeBD/uS8x9GCaXuEreZKpsciTZ/DHQB0xV0Q4r1NXgh8+2/bGYlOySxRfFEXqlST
Yn1x8QIPZE5up27ScHWc1izEc4iLxp/BrjV+n0GWyXY41QuvYVNOpNPtSlubg3AT
+uIMrFIFXaYh+/cQeoWVcktV7kfrLOALA52LWY7QJ4hv8qQQ+t5uns1mvTmoOHJj
SD91DwOEZKo1dCRrOErjENDH41ddg6YJldA6WkeFKk7ESkLD18uHyDL4dDAYCgxh
wIxma/5k3jzelR/+5jrUSG3VIVb/NirT2YLuuwaupOhTvm+YQqRczGEpddfOzzBo
Q98qq2hqOCsDJnAETSCRZdyrpbU0/9TAz6IScIwzTShS7IT7tcuNrR2QtW3CR8JT
2uijc8Eb8uu8c9hsd9IrDu4XJWWbX6FSQ/6b+yNuk0Y9+w+I4V1SqrhtRzb6FA56
Hc/tOjslnHlViG54jWMc6QO/CDY2iXid25ZZkPvD6tPu7dpIuZjjRMcY7ZxPkBJy
krx5wKr4so3lQevDKRrXtleCwiMtBNGzRjz6webskD6JVIZibQniYp/IKJ/YrELK
2wxraax+vopHVy3JrDdODTIsVs2PH0CCu8D/Elx8TptkVcDSO0AMWKZqFo6O80vk
PuxsCzdnU2H93aMVJ79AeXcNChHge7w7yHZh9Tf5wos5BajhDWbPxcuhHq93bhGA
a9htlRycajd9i8rImOgE5U0T+oqBcB/r//wpqEo4kshZoQnztdX12OFixkyfmP1Z
ukqbBDCTLPn5Z3v9IxaHQGHEZ3Mw5wygbXKlh0Vi6bO1BG39Kj4/t1Hd6kJ+bPgs
gBVlcZEcdHNEDFDtzyF75SdTL7HcZ1DxIEFSC25L54IYr9/VZw649r4EOpWcMMYV
xsFQ3wvpIRNkvtd7TYQ7VT/whxhnS3M1F4swvmCnO0QwpuYuayiVnjnvcqrVam4t
eFOtUn9EtalytjD/pHjYKEM0Quev+PMsbh229JEF8a0OoqRnb4/TKwPN4+DtMbl0
KhJ4Pt5uNa4lAM90gy9caIGCR6oF9KrmFCv0ULdcottgcsJAoZi/xOTd4TarLSmO
wrax7AuheFsqBDOjw1+6hnGyIWkOz9AR9yv9y7SDDs+kECc6d5ftV6RbKvIOb9Jt
yY0opPL5KsixaDluM7dbYZBr1ivTjaZfwifOasWa+tCBGiqIE33fowpOPOw/DhUK
EtuxQ8O6i8jjrOJQLagq7OE+LBnt2SD8hhRmTtMIthyuni3mvj5nWVM9xe+Bnty2
7G3MdqLGPeciL7rxxRJmTP5jlGanwoiqbIxGNj9GShNto8CVN8EGqxM3w1tlX+Ib
8KzQJi3pZIQZBcfJydHvyMVZH1/tjEiQkaLqohcrmZbUXNtQVVlOiYXO4KLNjkGk
A8Gq1Bm3W08D2m3m9EAwTwxHuc5eUPyIUuq976lBk0TFSGPW1vk2XDGzlmJHu9Zc
ykSgcB4pmYK3odIUQOhqkJPML/aZ3BGAviLGhLGGz03Rhfj2DohvTIS6LmPPr7kn
2lfycI+bcTGcP0PZFkQGsq3aCJ4u+wGRcoJ5E+bg4kfmJWsXt0hmpHl6MIMdVWf7
EHNScJ4dRPXJ/N6J73+hI7xoYFADmpMrlwWJlieFN1yhFPFFm3Lju91GyIUBby2X
yZhOgFpnjO8Z157GeVTXZQdMkMogRKl8DKcsRSp61fVj6p+MJr5Cdi1k5pB95j3Y
XsgutJeZ3TuYI34oAJZvycEoAtma2rhB1uESZjr7am31A/+gBgqRzEsOkGk+5xyd
p+WzuIjkRtnt0eFf203Brc5puDPrCHz4ppKDL2HDjBY/l8kLHCAJxhhx464eDGKf
6dV6NPQLHPvNPPr11nbYzZEdHa6qIyAmnJ76nTGT9wFvvYt9wyBtTRGJgwb0qmun
RqT8S/exgpJ5vY8dHCJjHEqib3Z5zO+Lx7poYAc+ttwGsk4G3nRi4sufC3J5yceM
a5QD81Kr+tQM+O2F+QPKh//7XKApyzil2kqSugxFOU2t5nhI3IOO99Gs/vbJtS1e
U4RVaOVQZAWXoWBlpumrOcUF7UyPh9Kjc/p71UNUsNi3UHu9lpGt0G5PmDb5P4Px
txYEEVLBrGT6P8fjLOM9BJlC5cwn8iqZEWyRXZ/Ou1HNwpIfDU/GE+Dga/K+HWi5
2jISDMZs3TAMeh/YCjTV9VpQ7t+t+tTJ7IXGFVIzCEY7zcgg18LWtIpuEQLrV6Ci
8IevGXjG84Hp48kt2Pdbnu1yvB+yf6ApoJiDWaqbMg0Rkir1G1TcObKMa/aGLCHd
HAGxkIRWHzdNZTxITxumw5wg9r3dat7z5DiBYHLh9nYsa7mypjMY424jX0afxlgQ
5u3o5je3Vp0RTMaeWY5F+wefWFRQCPmOOKx/7F47McwV0Ej34Q4VWBaIbmWn3U98
YtiUIJ5F0TGZN6yWQZNcH41aBYSH4NDXtHMxVDJ5Xfm30PIDYg8uk/RR2HnkXX/d
l6arpOOa3g4F2PIPGMm0X3D/PlN8JpUpKIL/11DRtZpnw8znK6yRPmzY0q/33dMU
hDmYiaM6sTyjj/0CRFyxYbJ2wuBC5FLy3JAXXDwCPit7PqP0b2/pSOlxB0c+fkmM
16Mj07pzp47AnvGb1uzMU/tEYkH2Fv2yKtTjRtkl2hAopGptzKBBjJs4EHXkulA1
JfQ5OxrXnm3xRJtXdXNCdFK5vLiZF0gVdQldn+ORmE6LRylFW9CP66C1ZgCc+Wik
+lPStBzcv+orsuuirjSJUUrnN8XIrw0W9PFaFXD9AUe0UwuTRWxlYsa7jV7oymoT
7FI2lbM17voQxpVbLYM/kOHsb4xhiGyf/AozmuDZiEiiXYdDbxeyp8zjSpNuzrrI
QiB0wt/WvhAVZEI/vR8OxPALp1oykjxOHxpB3c+PwI4qefZhxZC61TwcyNh6lmML
hGPYyo3FRxM7cUPbKSSXQaXbVzwf9QO3mIlzg/Kc4hu93GYK/OzrD9BDW7zQ/rrO
jRrd0ZSSKzty7vddY0fo3Vz1cXc/Sw0fScVLPWszaAxwnKSJdX0W6/KMTSH7KrOv
w1GJVPdMLxzehiQfSt/67or1PaMfTTZ0zoFlt/qfMLvW7WwPPgSpVg/1CHAmeGGA
/eMs4HUGijrtwiKquNyLGMcuH9S4NK/J5pZc6N/u0n4aWC8N1ommVW0sZsophs54
QAnzJmbV4Fn/xpQRi7ZJP15kZB7fygW6iIpjijp0PxvNlROckRkYJ6gu3FCsxA+A
Osr8l6vK8DGy3bUZy1liyz65kutxOiLxgaKwsHTTMLjk95Sb0QJmAXsFqDDh4OCD
BrG+xex3lWGrW5gt8t3SLtSvM80QqRLzYyeof6f05RGVhxw9Bz0ZD01lJixfGPNl
diDqdIchzVAore3udfq4i/xZ3kYrX8D4mqT1HU5CDth5SXrL/LtEdhBRFaoqL9d+
ZsmWHwdj+9pP8PKN5htohDzKp99trY7IPv3d9AispppAu5dZMyDWJ8ogeoX+IjLL
fxXSEYIosZviqLK20N8uLyms8IdKRG84GKNjctTc7fRYBEYzTdMzTq2rMLApfy7M
9GAAz+juWUWY1VLed5nwF6Kr+d2eLH2bvBkrN1Lq2/wOld/FGckcSxC2YFqoqdfW
RDmUbyR2Vr6avkEKOoSXS5KJ1PMZCFj2Cg8khs8x2LDBVUB1JaV8S+5KGWoDqyYE
Dk/rWpb5nnVr5kYsBWmFazqFM57HPGyNd1ULjjsVNvbLec+tXL5rPCtnsNrn3JBD
bcXy6Ts58QbgGxZCEnsH0XWjVobe07jAK+2lY9lyF7se4mTJNeSszYTXTzQVVTM3
MIYIm0HevqXQdJp/Zp9JYtI+6tWRhq3aM6AjNSU1W3uzFScIuHb/jiYSQH9dmYKP
JfxIEI7W9g6dky7jTdsJBBWeWtDYnXZTBA/H/vjRDAiPEVQy7FSuYZyomy1KfI/V
sC54zbGfBno7ajOzXxY5wogoBwmTxGcRgb2JilGTGbN6Ivz24sFtVBGTgvKjhxsK
oOCrZyclbKXigucqE9lW9zierkRI8Tss2dUGIR1/3q205cjs6v+mLaIGE8JIwk9E
OaFs8tFG8OJFyoUdoyZokFH/bybw062jgeqt45uA3PUMDZHeSKqv7ntbTaUULwzn
H6znjrEdxtNpei2AXUNa/q2rqI11rBvt5P6nThYR4ExeN7sWCeWS1QcWX0xqSMCV
qcNsDRigssLJ87qDjhzBDx04mzXxSJAfL6YbW2TIvSdQTDdfKYzJLNSZSjTIO6sN
/sJEqAfnKU5RHxYSxOTNA4o+SxQvYzmZRVgYWos5sYhwIip3azMqsykkdM95CKtn
Dg+FGPwoUmv242dkvKCG2jiz/8mi+AbgpMSmmBhBUmLEWwZ783MUE84Y4mQ1zHcZ
X62aLGuBJh9Zb+LxrVWNglogjoCL3lli1P3OYFHFJG5bATTAra5vsTFS5w2+LtOk
LqVKG3HdjR/7B6xzuN/q3zr016hENIEvJiexr3OXXulIl+y4h5Pqqh+UsxajXCxw
jqFtWIOcVjF84gUsUcqdTK8vKXdeGLvvjXduNq6KxWMC1AIk2REr15nacxgY1IX3
Zrzl3ArHmdAQ9ogo7TvMCe4sKtPYqJ1rpEzVhglGIoRQwV5Xp30QeI8n2VSBbO4I
xgodh0oKEhoUQalLuX4FCj0ZgJndISq8JX+NMJwhXoNvuitE1XACqKcywp9ig4ut
BYHAC5OvUwHsL5NdXqodLoJcJOKGOUDhsuzW1g9vFSuEX1tBXrgqKP4VCptZuJta
dfOvKOMfBqqPsM7Cgzgztl3axdd1Fa8n7fKcjpfEua7+KNs9OPG89hvftVb+sZw2
X7kguybVvhQY0xD5/ccfe/y9ogON/3EZAKzVp37kafvdDEeCgdOsTimFy/iRua3U
QHdHRklGvW0+vRmlIrDKHDzuLKyiU1LHmrxnttEjVz/frRkZdo7SgWLMtzOdAjPe
0BtynpMezTSfF5Dt9yTxTCMq/3QmfMBDbV/JxCbaPzLrXrTPnv5LZgTL7ZUGdWnC
8j3nmnxBJVNGyo6Duy9dVXGXgMQxE/uQpDnQZfHNpZY80lJfUkcRUovPIijNhk60
JoH3T8JmsiP3oupdTtUQjHXJ6/OavfAuDX/sGRjVgM/wQaTTPI8IOEbWzOWti7Z/
oe8Sx/OKNIf97b2nwXX/Bil0Pl4KsgbcPOFjygnFMNOJPl38sEZdCQhs59kyR/G0
DTlt3mRHdfi0p7FQLZ1LBwja+kHzS6rr4sOOpDiRYjcJfac/SY/n8fGv9O4w/q3r
eBEle+SCbRnGndwdW8qY08NnY4AvW2UyeLSyebnxSikaTmueY6jar+s0PZX+sVo4
Tu+Tg6gYJIPLHbWRcX2erk7eprsYObyXpxCWa/DuOZuSh7AfKAOc13MgYpYK9xYg
AmrZGG1vvycWbVn+iRi9GK6XIjUliF3dYrKcCO8KpgZorVTz7JUZjZQX9LwAEEri
nBwnDhNa8M0YMOYKdHVF2mEw6S9mr7Sh05WbxF6Rg+YBQxInUumvaly/uvDT4UKo
yglVZ72aWlyy9f71PJWGjlEdIFgz0f2RCtni6O4uYp0hLwYRGmWVRidn4Tbw0Zd0
3Mae6L5eZUFuj45TNH/5s0ttWnTy/crZX1ELwTWxuAde54c+sdMTGZ2k0OgL4iTm
AI9ankLc1GtWi/ztYUsl/oyFNjisv26N7ZfStiS5ul08/Vrce2IAcm4TUCIq4XWF
rPg5SXBo3ZaQHRJ6WlOW154vcGK8ezCtZfBfM/+gjc29UYj78T9S1mJ02kT8cr2p
LOs76PRJFzC115Uoil6IC7aD1SPmVW6gzncbGAP/atk9zXpftr3p1kmgWUMyTOwP
q4D+kpNpbgv45bglcfqfuuUgejqrk7SxaRgCCfoGSBZc+L1SfqadWQpe/Ztw5oVv
so8+RufrZrmKhQr5YPO3gpixtPALr1yyhA5tZY1rc8G1GEbJQjHJB5auDwT+IDJ2
odS0B/YXOkU+rw1SySUBHN03hPFgFCTZUudaMsbDgdrRHaKY86qtHRzgf1eRx3li
IP9MfstmNhHlrvnxrNI+S07fS3i6iSMORqbQKod18alU57BibtGceA0/bugbT3lo
Ot6hFeUo1RUNXlQZ3k0NITICQm9Mkr39D/yZKKglkLv5IlfobpypkXTlICbetfsv
icTWtqHQ4tLrSNYjzxqlRNSZsJHGP9luhdIgLHV6zdMqaa9cKze7AL2ab7lif14d
BfHhMxesSDvqxiJ0BMs944VvEwPiESa/ceToJBgOjnNOpWZ8FaQ5KSzy19vr/6yf
2Ksvkr8UvZpP9rLWZE9qzZh1XrkhHlLhIpYzN+09Fsu14TkQrSHg1LvYecMk7gR6
8BSlqffLGvB/eJDc/UiOdO2Z8BgGmjG5PVQWb1QWQ3GsPZTv3Q9BzJ9nExkFcEwi
iysGXFXfwntrvY3FWcxRXGpaEMGI2Jc9i3wlvi35IXQzQtGdJlj4UBtKja3I+2L6
K/wmnO1EU4q8m8Ty2mJY//kyxGZGFzGcRkM5QvCF7ryQBIFo4cQTrYtmeR2RyYWY
hQyPAEmxBLvWBKb6ye2VsjQ2x557YO9XghWgRO6Jk9LHQCl/Ep3LECwtS0+0P0LX
P6fwIKwT9YmYj82eDC+/LH6n4X6k6WRnvvxikbczMBiUybdvwhoqHJ54lIraFt0T
1vmVR/09SwgwMQ3h4ZT+9qfs3SshMaUksQRzzgK6sp7YAJ0VPuD9aMdIQNofwclZ
HcRy50VJ5Ruk2UsFu604RJoGzH05nlAOwPSzHnewkyo5Zhx7FccWxMFo6PmWXc6e
fExU7TJlDD1MBSDBsMr0oMnpt9lWJCaR7y1brvXS+hFwMfYcNoTD00wG5ALScYz0
YXAtfKKc2kv+VApEacuoIzijDnJi08Xe9Wpj33VLSVtB0nSjV7r3Nl1JjM/M3ttY
FXyR5c6I4N+4isb6Wx4jQD+Bq5i8X9gFU6h1R01AhH/78kl6XH9X4VeHArNb4+9N
fSALRm6nPMHWZ5ReatearukmTEcN1VqrqnkmXgnd3euwrwtA9zUaxFcisFkeEASB
mugcOoH2hEGEqin/hdt3hTJ40vxLsQdSnabg2CWnCM4TC7mqVCYiYg1l3X4iXknp
+NQhIV8uCtHnA18hFSTCXtE3MkHSVrm+BQ4guFN5dhm1tRmpB0CKJ1/HBpgdLoUq
6wBLdVR/vc8CJ73vKDb8adbqbm7uGAM67/qcvxyYLCCCA+wS3gPl/rIcLWK9scrk
YD3BpUJAYdUbt8l+KGQKAOHbMzpyNLHC+U4kcMX0QSLXMRaIsU+F+fIEcT+gH5Oj
rHSgLN9mruRO7YqJr7H3QYfGrgOMAuFwCaqp/GxHRUiusyMKPJVjAHEltLTM8vGm
yYGKST9dAVps4R0XaGVejAdcWOOZlBODKuK5Gyb955LOVuJmQz37pX679WewzZTu
Smc98eFIZvMBrXMgkcShic+5zylE6O/dEx/bvu3HOLHkqhtF2mVz2bjEIlySCyR2
r6MkLfCr/9pqwe+7XAcmQvuWFueY9FHKsEODgxwDuTX43BeYPIdj1UM5jWOcl+XB
n1GTzh2xgvuxAY7QFRn5z+zxyNvn6iEr40u9zVXdg0/RRVRRk1zmPk9pCDx7SZtO
EhNS9SGnoUzz1KbcYXxkS+/3LOuKwGqfBajO+jbEY/bceTxBM21o+XMWU0ALqQba
mW0MKsw03P3T+ZmvBDdfR8wrnLKmQKqugdG3H+Gig3eB119KmCbWIQqStFIVhB/Z
X/nRscxuygcUk6iXb+9HXgl085u07VqU+Xpn8DEWSnvqV2WhxhiMVyhHWidYTmos
Z+obks4EMjBSOcb3QkjcEdleELx+0nCkJX0J9EPLxKyrL4QmeDX1plm0hvQrGH/F
6qmGIt1hN2poCtL7pyajr13ubdFvQSOJqSollwG7TbrtvSuB/3mFmaQOwStDRPBC
S1q4Eko6kUCzh/jAKyFkCcaJ0Nm+9VY/laaIgjLxKn401/UKs53Car9wYiLuYYG7
2yLMLgcqaLkm/sH5heZDWSfaVpLbfzVnXgJonorf9Ex1Ko76vTLAjCdtdO5kcuO4
SmHgOYt25c0TKx0pETS/s1wmAExgg9ByTgOQucsYwWgmfcqxbsbqnI4lcYjisgFn
ixYGT/ZQjwGk6Y06FEmEIgMIq+t6eBF49YOgOACpqsY20j3m64lhjOOhzU4IXqo/
d00UAupeIbXA8gi7tKHoaREMyJdAv1Pwmw+ZijIFqirKwBOUvXdBbugPKXNTSSdW
JF+MF5N4Jv7k96iP/TEDcG0zS7nX/AgVO37kG0ZZRdGKbzLrt22quhFn5RkC7J7O
kvdXvQ6HE4Xwkfvv1Ww1pQ==
`pragma protect end_protected
