package avalon_mm_dcom_registers_pkg is
	
end package avalon_mm_dcom_registers_pkg;

package body avalon_mm_dcom_registers_pkg is
	
end package body avalon_mm_dcom_registers_pkg;
