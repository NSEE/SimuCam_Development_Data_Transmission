// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:49 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dWFux1gweN3YJlWiCkvCR3O/PaLMbULZyOo887BVE1DCpVMcxtiFBXu4OAC832QY
y30Yk4IF2H/KoY9CVeghCwgpExotalk8hBcb1Xn3xomT8mqtjg6rx+1PbKkJKJEe
yJVQSyPDEe9eRUTetQDEsiG8mSTvZ6X+05uL6W5tS2w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 84960)
PqmrLYfGMJDxyLOCXFkkUcD6r2AevBj6TSmY+QZKlSmW+eU6GuiN4vZ07Cyb988e
YYV2nvcBnDCgjJXahBsoxkFrgH5BtdO/eZOS+dr7tfhHxwaUIXUZzpeegQOO8Pmo
QAm5GZI+ktNXAx79kFvtFQ1BcAr/UAenlb0TZEA46afzmrh1ib7UVlHk8JwX95rm
Qez1/UAcpTpRUK6Vz7x2x7iB95vfY2Z0RTWsONIZfOs3gKTvaa/P8XCq85jNGhLt
TYtXccJJ9lSGU3bmE24Qm3Vipzvdmc8WHvsNv+xMtk7htQ2tXlLagUOw+41xEbH1
EOl2pYZws1p3RHZh+kZLJH6CfEQVmm6Cw/w1MIDhsg8WC4oXzuaXsdPEIt7IFbFK
5cgTP/DmZW+rzaDPTWi2koN24Wxr0rLuF5zmRNvO5MKgxni+w7w4fQE/TKWqQDv9
NihTu42Hq36sUo/8DsOFF9FB4rx25CFCC7lmKehPknjkBOGF4EzXUOvnXNrzRHK+
7wQHoS1f9r3rsKW1FMdpRfh1XQhk0Qo9lk/vFSPk8pYzGAT/REmAgNFDNJjPcWN+
k6OCJX9Pd03Amn4AC2zf7d+zNbmJQlUPxfB75kRkIUMuXNyq6XDK60pD/SQ8lZ5K
d7o2BQgFwYdVFnFfTt74650U6ARl1n5Oc0r9r8hMRYeb7dDrgSwN+hKObf8bDJH/
7kdlFTc3VO6n2qh9DpweE8EeZ8nubeQrtzhPvXK69srzzA0WwGvIemEMR7dTN+uZ
qUPB2Ejx/EUoPqLXWixxiw+P64tCjwizwlOqFGMUoSpcJC/DRnLBPxVgbPAfDgHR
k+kF7qCaCHTM2K76pB6TnaSk0zmw5GrSN4vD/rT0BsmxnUNzX/fmeB95Drw3Fd0l
SgH/t3KbM2DZ1+E/zRF9w48V3uXKsnudzTRRqz60fjo/5KOMZkOZ/Ag2Gu4LkEPE
4tZlcmawfbclg8FaXjfxNzdn/ibMrFASqtXCEp65BpEnjf5LuDaeuBJq8t7WwBk9
R7gfQbkws6qafi8cRmhYdaZW2t0nnzvG3RdCW7FAOu8xe2+0t3VyGCY4Egj2JVkX
k0LKJyhRPo7gH7IQAOYWrhTnJVFLQxsMDyc8+v2FA5H0DzhYxXyNqjFWino0vhDb
UZmSQOYtXC+1n8HTsTO5qmOZ32GwEY95aklTkcqbGgAaqB8PPaTOxk84czk7oKiK
HuPGP9Y8SH8/6/m+PeKiXpcSePOGXsT3+y66fWMsGrA+LYf0t+YPTDLwMTVYKKnL
ozOehiCtaWuxbqixtNAvUCv2tnCck38qn4TSnMeo03pJ0uPyK8re5v0pdH9T2kMC
mB0KIvzx56lssRzYlfwl4TzDQRIAL8C8+aJ7dNBCQppwmfnNqn8zo8qWFh3D6K06
Y5z/XnJkgE85I2em/GE0SWvnha1opCOXomZCKp7R74j9FpMFDcWMgzR+ZTboBI+s
Xyp9rXGp023z/NPSWE6xMk5oUKV/b2gDOw2DXY9XjhRJR4bYKNj5NFk5o9LD3DgJ
XFgIe0ENfth9/Kvxka+D3bsaaAUDHr3AFe4kcJOm7aQ6T9QMc7AZZnFTuBUFzdoT
DLZLhQpYvrmPiqPIEMtD6ZpAuMxDj1ocF8UQ/Kj7G18pb2g5GbRnzP0Tpm9rbnbm
16guanF+CPUW0942jpEdM27b+9kyfhSZDjtjOVqJ/5mY9pEmjrjFp+b3WID3Lt0C
bEvj+PuOVGhUryx0m2RgysTorsjBSvn48e2RbTQyltXvnZ5dL7sDN6yh+BEuVvSh
L7VutW6txoISpfZKYKtq++No4VM5V0x8J2h5NieJJWfy9eYhiZ3wdXqnNcY/wgdB
aAxClJtuB7SS32DzwdptfxJChE8DtDH+nZRFy0+mKVTpPBwKMObCEtRt6lh1R47x
d6/WB7DnxzuWlMNFFLjBxIw0jon/32AlLQcERjOdkQ6bYePdlWg+QKwpaddbXzoQ
X0VStV33gSOiwPUelT3yvlyhYjhJQ9v/+9CxdfpAH0Kf5goLXgqpu6bHK7wG3XWc
v8jOznGDxa897MM0OEJStY/Ax7zksGwIJt/sSiVTDjkzWNv0pWvidMdbt75HPRdw
MM9XcUj2hdib+G/rKFNEv/aK3YN/itnQi1Oq9vDnf3I/pb7h146UNbct0lThpmif
OnNI9hrHPKHxfATLO0xisjPvM79qs04DGylbrOAVcWu5L+zKmqU7J9sGbBsRjWYs
Pbeve5JfLq75B9Mpc2/Nfj4tIckNn60effpEpNrdDIV3WB4pxu8+0zYxUHwokz2N
eSld42dkAn8DQCTEpdl8qUrDIhysdp0n9vQsbhxkd2QnXqlp601wDJ/Jl5c2uedE
6xBZnoJQ1Pqkpo2deuI2zKIIJpj/UgphHwgow4rMKrdsXcYNFWb984WKHX7V3ioR
TYPQ02bmMx0kIVTeffmonAwvpWnYLI9HiAXPYtES0ErC1ZNOjdAUzTwXo4q+qGST
Ig8nuBi6nB5U7DZN3i05WUYeH+Z+AXjI/a9GRwsPR9ZGfz5wTShFDDTq05ysphsT
0NTwjHeBHI6QAzEQVewwJegdTa61aRP6w3vTPqAuxV/WeTuwiYglrB+/VFvTF7AH
IxWWvAYRYUs1TvWQLph3RG8o7Bu85USGWvCsaxb5vX3lJkK+pLPSmBrA0mrmpxyo
Rlzd4Rb6a/IuWLmCwHyRwpc22teBH5gFKHB5SNXXQMBU1w5KseeczzAUDurkVI7d
WUc5ZjMLmMy3SicQYvw0J2+x4kJcemTlmuJ7pq89u04cDS3iQjWSD/buXcPCm2lC
htFLevps3jC/34fTnCvAC3J/jNRTQw7upHriq127pvfk0qcV0aA/PrGqeNXJrPjA
PxR1becKMkBzXrRad5+Z6RAMFy5uiHuFb9qrgbdsmyTMk5CV7YelWuVXnmoLz67+
WWVqbMzaH+m+TyVkFWVhvuDIJ9FLIkfpMPPPHoyWN3HBHr5kB9WZrJejNjH9uPzz
mGYD1ajPIi+1Qcwg2/DP/MmL4UZmg71Drw4WMUAHju+SpMGvH2iZlf9dah83MW2J
W8zo9WKQULKHVZW96nAjarig5hMlhHokPabMMUx4ckx86TTnusZES38aHnC+wuR2
3B/8aebVbcfupWV2EiXtJe9FjZ3Xg6fKdfaXAWm/4Nh7Euwbefrek7CPZdXgdwxC
PtN26E1qEMKhnZTk/NP406aPQfjQfOeOBdHAnBW34TnAR1HqhUVVME/2XYFwuLZc
blhs8qRQL4h6jXt7lZjEzG4j/QRw3GtbkjDsXnCo0nFhtwyI2t3X+bRs5bWa63Gy
zEsXHQ34952n4v4v/+6lujky1LSc5Yyxv+bzVTS/SLxewOuztTC5quW5ick0gTqy
Rcb/SOMZbtthfHyELmeDKauSbavDKolbeG/2LSKvLIxj9QHslzxV/t6vY78vOFdt
mGqhC8XkT/1NWreXd5MMeFwGZM7LgrGeySukmsRT7trxg1inseqe61dgwZpsWY2g
TiBqx5hptbJKYLF1lLG80Ua5t2Ot8vIBJ+4V1niojwhm4p7RyKWdqrBtSAt6O+1j
d3nQodBX9Kr7BOqQlQqXcJ8Yek3+jjWbY4UuJ/vgu1xHCC4DHJy8W+U98zq40SWn
LKWAmWeqsrKdn6Y2V3DVcQ6c4N1YIGZcSPL01WSHqrbg8ZGsrNLDLaMGeND4lxHp
RGuQvCR6Yco7lWkR/H45J1AFR+NmvDn8kPF0WAoRlwVjNsUWuTYbyuZjxyNYgNg4
UNlBMfWBYaqFmv9lViFwPMxe7JjO1eRxngutCG3T5D6LcKY9dyfFWtyJyPXIoPHp
TQUDnw7CrDfE5/xUNlv7Qf24hFjvdRrdaSnrmX7s/pNok5OiTGEByyHuFTGFoxph
fk7OS+3f6C9VzasYNWgUECUJatvoOGGjtGcwyoDtmbhayuh1LVGLOeRxqsOLnAht
7EShs06HrMnvzTkxxag56QSpCJkzv9LKfD54+LWGS2FjotQgZUwUrmnKMj5FfjOS
OjeH8AC23hzhi9lgDagjW3gYKondERDEAjOlv7++zqsuRCdQEU5EFPIdWMs/tT2x
Lve49D23jRz0k4rG3YhepKrvQRVtICQdAYzYgt3OX6s1Io84plLx1GgRHMNJ/Hb7
MW1I+JxX62OZWTFWGdW2hcof3OPY9pzyT/cz5W0eZ0CQS4OTzkQVGaGujtS1ZH/H
Px/0l7W9gBfd7yj7t3nJ6zEi6aE6Cl3wouAuU2WmqYiol3xZ2XHzL6ClWroKwLK1
GBfMaSxC55uEG+bDU115YZwnG1mJB/mDkku+gGfNOSCTsGbb4GFSiDjJPktTLieT
UlBaR5+HlvJqFpOi9DRL4ReGQGV2Mb5FbDHRD3r2kB7xxjzI1XjCcpDNCO91nqCh
JeDLC1mHSntSLz9LCo564gQBxllJqA6/ICZ4C2Z8Gyd+YmBY1jDKO8KAAE9Gi8a2
p6+ZS19DREAH9FNqvHrDdFc9OUhcOKc6GZgq5tqsLfC2EQwaQMYTVI15gOJOE5fa
vOGiN8Xu8yetQFTuC7zAAcOWjUUkl3eFTTJuSRAOkqTYMzgbvJTRpHtE6tJivx95
xxrvG9T4dx7pr5+uhqT/cU4n5Rg4Jef9e8j/N5AGGNUbF+IvkCBm/wa4HPTHUqK2
A5elb7uexaWJHhRj5alN/53dc9h/deUsakDj+L1vVAMimAB+qTlVrB3ZYTIFKmzp
aH82zXPEfg42pwT2//ME2FeJdAAUB4/MnCRYIOxrsAotjQAIwJZPFDEB+rNg6w2s
3n1ATccnabsiG8mDzutIaVIJASfwsT6XC0ECafTGhN7lY+F+ph5rgyDrN1GS3FkE
0OLXAAdZtQ7d2apKcoKl7SM+dMiqs8QKaFZa3hd00W6B0rZdmYzqBTaeg6Kyg6lG
8DPEdcIrP+QBbtr7XzcydfUWw29yCoR0lj+365A0pH84z5qklaR+F14REs9QNANS
t/0Uxe7IfkY3XYzfQc4wusCvthMlzdSWthUtUFSOU5gRG0QH/CmNVHeA6RIXYxm5
AdeLrdgTuuPilATDLu+r0+aIbnGt9N3PNQikXsAoymtrFA0KeLLCZjOhvovyNFFS
ohkZL0DtEPCiVmUX0eVkuhRpwUijfKLbppmo5jGJsdyFb7x4zR9jmwY/w8UMeFub
dx8llMMPcNKqBxuAPXWfogwlTL3NoG3vKxPLDuML0d/u4fkdUUpAkUZP7B3iQHK2
OUA36bV+r6shEjj8nTKUEy5okK35qI7u+ONlABlvcvr6DIsBZrS9BUGLB8NXbfMX
yTIIM+s4L4pnVST3pM2BvQ63TdQ02V3FqPFgfb9t7PMU9V61jtQgOV5AF7o9+KgP
BCrLUTwL13aKZTxRbHiGJem0buARxlGAq2fKHW77ocR69+Vvjk1pJvVAcjbCwqoh
atX46meAPBUayViJj3RIBQ8oVB+z2f/KsGRmiGMqgKuzTW7yDC87UCGuEH5khXYM
lPxZN+WK7cWP40znp2dIOR1WYvHBI1KdCXi4/vSpgf6+qjknSHNUHIWNNFBHqjNr
b5PFsRKw48crIVVNKvex42l/sWN67bcZzXC85NihzqQ4Fwy6UNYa7Wgzr3po1U9H
p82k++VYwwqUFKq2GqJVNZhptc3/wREOwgiVW8iHRLxNy3GjVD5qq7B2DBpw1/bW
hewh7DVMQh4DRqJYwHk+6qy1JRRZhW9DEB6V4ap4afI36ULhaBT8hVAaG+dA7vIU
FQ5OnBAzUm6PN3usjasix289H8anB4WKpEorBFDL+R1Adqa4VJwfimt2+OkcHi8F
G8OhkE/gJSpqGegXAGPgDuRkB3SL04hUBA45Q+S+UiiWsUugnRg/Lhiw/muS3DLs
E6Mc1zhdEddsG7aQS0P5hoBlxRdq/Y/yU1PI+1cWfBEM+EnI7NLlAqQ+idy8Anql
c5FoZwOaYSK/NgB++f8W9CCNcMzCWkPm0ac5VcDgVzb6WQTz/GYq36AgrAVunWmU
ei1lw3wZjU/1uDUD2DD/P/KHFIpiaEHyHuMgCXLNroVXInfZywMjg4bGFfkjA1mF
+XIVJH6GV8HtWeFTGL+acitMiRQFovuZoWihwpi38sQx/LQPBZDlw+NDU6sdV8I9
9ZetimGTOfHGgFXuAh0CoKlgxENAscRoVoaejIggsXhVEH+lYlDFV4/NdgS5xPAM
GTX27ncI62JuenAiA4w/0jcyvXaLGWg5vuWkOgBU9ogSJUGcTUTcsrtvRzzwb8Ed
jXyNdktzLwJWmpVYgno9yb3ZYUnSvAtIDUOvzC8A0GOmLjbATRc4wNxu70xtaMwL
eya6cA/0llf/MkVXvGw8oGVtgWjkzNSHWqwDrh9+9wbiG9Y5kNTwD+bPfNPP3wvG
EuoenSWMyQ+fowL4p2+2yE/XoEfq0/UDjrGtSpX/6bk6ctLCPzqEdt760DYdbTUU
ihtWKC9KuJ/tMrMxr9/lrqAFp8TTjIdg2rx9PBTTD+6VvLt5pACMpdYNvwcW12H6
AlCWZYFErPLDMfDhNgWQRBaOVKutnwWi7K/hDdUSXQ0ahfnrssgVh8HP78k8SevE
QIJgZIONgVJeF4WT4cB0raf6182qxctUjrWxbCkmMJjzmsjE3G1+GKKO5rv7yRrY
7t4Z0oOfjBf8hdG+e02hHFlRw/XI+br6XPo7hxHtUbooptgo2kX2j36mMxEowzQf
VJhIGbkcJYzJpGnMdeFkaBmiPaL4sul9FsEoKbKa9Hpx0eoXcKeMCv24I197OLw0
lIydxmhSfvANlBphTwsno1a84YKHiJMvtapj6ZVrj+VtUjb5HiVlJv4Z8T/TyHNN
uiUlt2x6UE1/cN8KsCoBll4OGM8tbQB8Cp5GQ3SsLSfLGByyKxwhJHn94KvermVv
F+WwmvNjuyxdmsU8p0XC5Z/+/d6MzhZ7gnWL6mcVRCG+g7H3sJJofqjdCHoyOt5z
ycecPNKYPkIYIEuvpoyJJ2pFCsWO9qyiQ3skDqTKzrSUXD0UC7bdnrQw9b1cnlKs
GSmZyUDLompXoo9en6L95HFqEuhz0NJqcimiabvrxOdn4OqyX400UPGTpEKHR5gF
B/1ZjRDo5lUwPbWm0gitP4DXswyFCL6upimVScszcjIc7IrzNlFnOb3tW/x4FYdZ
En+M76pW+D1r0AOlGZgV6lp6ccYBafnnogpAWF5jFqYGhDhhg0ALX3sfLUAUt1+2
rUWn2eGrBbrkCsdKnufD8vVgjBcSpaIYpynHM0SAFe94AFml+V7qjx5905QLB/jL
n03PqKt6V29FzjUffQzhFMTJkQ/6Hv2ACmGCriYeU2/f/PLo4qKn8V5vTlR1qEzu
KLACl0lxZqr/rAcLYi4jNZwZSE397MwPzQvCUKaHLblMj9DlvolXm4onWlh17yFb
lwNlq3VG2daiZSVbARRxuUmxuNpBKtWhA0ifCdjdFMOy3hCHDUzuAx9diq/Cm44q
oxAIfCy2AGcW0ugp4MmRpqBHjJaCUAzrgj7bA22F1N2RpXv5bt25XvIfWKIlS9aH
t7hdh6xZ4nWtu1c8zKpvjFoK1a7FCp0WDPO/+pwBlYBKuqc2pCHY6hMFI6mxY+Wh
aQx1wdCsndmBydYpFn76ceDNr7cHQJYZBBMrIO10l0eD3LL+3EgH5dBiahryN+7J
Hh34ANjrHnX93vBYlUnrifcjPDEdA+IGlLMvTRkRhBN+kINmbshSa63+zNwYCTnk
q1wYkQ1lJI8snUKKFspjQUJYJpTpRoRCqzr+UqBUFHueCYR3WqMKwZWZDh9m0DQo
NeOxCu2RloLKKdyu0+Oe2bIuHg1830aTsp+NBRimVvqWGE/UJKkryIYKoKix/7mh
t5vPa7Hs2kpFXzpHnq0ZVC90gKY/88bVnfNpZszeoxvbRtt79CujK9NWSsqQB6Kg
3MogeCs83XhND0SP/DkSd2sTPodMDR0ta5XN1jImmNscm8AEhBsBKMhKPac5YPgp
uK+nQzWVacbULSdNRrwdXYY+zXpjoVyCnjkbMBj7C9KV7+FZLnG9IBgCJBz85yK+
KkM85bkjFmEkjPL+XqlS+um3h0vEpwQEUM7r8pO1qc6XwKVUJ8X3i0UUDxVzRrAM
WtieqjIJQFH2noBW0pazdRJh3b9P9UbhrtXZrXy9M6+Cs093rBzsajI/MLEMxjhY
Ry+RlnWWzVUOgjJytJ1z73lKKy/1UM1+YTm/swiNjCzXbGVHNoSIsU3CtTm5ACYQ
Du+8Qt95D/w2hDxfJ5OE2oUNnwrjosLMelsGf3cq197RfzVnzBV72jsSJHiwJYr2
4/aQq1/ZKznOBnxLYcdxUJ/a68zSkcYR1i8NMlMZOa+GRcQjF448xgoo+NOdcrkP
xSS1rpsOvMzly1jSQ4oP6teRu6Jjt6+wkwd8pb/7clkmg4Zj/R6wKycJuucYWICj
2a4BtXx/lO6Chy5Mtx90C3qMYdaOOclOS4xK9natNgWv2IPUVFRP6tSJThBmQ3Sd
SBmvbyFVTS2gsx2ybQrD5uSwPZ93mZgLDIZAt+/9+X03lVOlmFv2OmUj0wFz0rYb
06OUE/fK9SNevLmwT9nhhHRnjPKPnFwJFS7agp1JRZvooKKQXYi38/Ff2q3y2bOI
QvGbiw0LYEIYs4l0r9IJuqUnatDFVuYWDlszJhANIH0NP+J+D8NVes3sTP6LHlBh
pPxL1IKuxEymsyClcYro+mmE1AFYpqJ50RmeoNn+4VKBKU1tfAzU0/rsV+XlOAde
tq1Gf613m94ZDwv3YzT8VaG7WjJb+OiMxtTtn0k5AzUpnY/olsyCkJ/Shg+ZHLsg
rRHFDZR9j3TMBmP96Or2icFYro3eog6C1zkkDLbLQYCgjGOwsLI+2j1cesAN5EIf
YGDVrC81C/axz4HfYYx768PwrpxI3PZssfeGEE0k0T1+q2U2YGvwLaIeJ4SIyvn7
B4H/BxlFS526b+aenaGERZTvr1TLMNBnR1jx5Pely8ncXMRyTeD6adYHaDKpUPUS
8alfG3Vj31XaDKkT7SDB4QahA1vEQBhXrFK6dlG4wM0BqFDuwikSxHcG/Aoxx2Pv
raVUI7ZBG4Vx2iY/BC/l5TGgLWFNLhi/NIZWgd+NW7avq8w0qCorH46jXm+RQ0vX
ef08dCQV1wW1XaJsnGHq7bQNXGRfOd7L0EAGgXQb2GSOrHO9ZHcka7w9/zHX8y5b
rLOkp63G2nOTAAOriKH4DjQV0j9NO/t9eBQ9QtnS8B5w43uvMF0ZeCfhsTJh2eCH
FvGCb9qqUho2LTxRy4t+e30P4n7dtBjb025uQnP9OEPscU5q0oc9unKUH2QBoHbV
3YdU65lzH3f0MJj8T7egjVlRvvmo3r6VfgUd+doJWozv1IK2aVSblFOX/k/3TTS+
Kdo4obM79aieEKLqs406gBjlFnOieNxVqi2gV93mUf5ecG04qBOKjysg0InBEQ7U
BfdKF4X9XurDOtQeYpe7zTGE50L+K3knFe3seQV9ES2zs/9V5Xt3OUYSy2nwO4vh
vayAiBM8ItRUbciOkeWAFzVDpUQSc1d65sMWaN4zr79NgXnpDx7hqisFvV4fdELY
UDs8HnwvXkzkuFA9bFzyU14ss/J5YH06ojy+kneD8jiK1EOXH9KnjBXVX8GlSTtM
D0SLq3sGi+mjHTTM83e5STLeCKJo1uSFZDQsBGidCpk021h6FLGPC6PCQbHhIRxP
DUDA4e+d5E+faRcr9nLtoBoWU9S4pmzDQQ1w0MWWO9JXqOkzDdoz63You4tTWvoH
Us2h1ClpfAtmxqpDaREAF4iWXjgGItdYXKL/E5TZgjSB6locxDqE0pD6zv+eVFHg
qui5hF/PmaoLgntVP8V9p0daSkEFnI3DoLDtYaGVjPphOpcZRgbLBPdX575rkdzT
g4fthnRHYypU2CMq+TbPBquBYELIhaFN477cmcmI2oq6dR7VDe4azfs9ipWjIz8+
atX4afFU75bJL6WHbSb7F/WW1OY00PEYcUF0bnWojnTQeMgl+andpyqu1xMwYJ5a
tJ3aO11ez/xvdTmHFQDk2ErXZHyy2dal95dZ/2oFhFDO68nuPc9E/VhNzyQ/dvEU
ytBLilmHZ4cb0nmu+fDKAbnTeoS0mhPgYgpE8BDDqcTYHfuXwPTeJD9WfSGz1/U1
1YVQ+Nk62meGA19e5yeBE7vmrMhbnLh/WncKXgDGbfQsXHxOZjlYTzSW6vn6hB3h
r4NerLw0ba2ZuV5kaz431yHFGq+Tzc2l2DdsF/XpueOshEpn/B0ISIr1eOSe8uXI
LgtXH+rz1n6FihS8tXYOl5GXJZFnVBxpfhHHXaEe/35w98MBDXy2zaZ44rwt4RRU
rathY1HHX+OpZdBAOrgsbLB1UH9sA5A2RkfsWmMavUM6OhFhKZ/AWFtwnDrsQnTU
JLYLtmbaUPdyJ1ReP1O+79OkNzR7jxZmFFJXlmtfMvukRCulMs+ZkkcKuXVn3gIR
zCSy51it1OhNEHqX6sTryyX+wx3LpaNr+rIuXb9XWwl19do6Yt5X175/1Wa3XK3n
yjBQzbY2utYuwzNOYm28gDNtVJ0ng9sVh4SCU93g1mBi4A3e8lmxv1nA3lpV0ttX
0b0QaCqFXi/+G+49Q0uAWY5hy+ex9CMFmOmp09WRzEXndwo1ciFxe09HCCH+o0xc
PZ6W++d9sa+vwwiOov983dScqBdkhIBK4ETNjeB5aKnUUYLYbgXvEOoeP0BApTqr
MXkempvZc39ohnjbxueY2US+Yw2Bu7ZbB0uhPO3a1LjpK/IztZ+RGcFSADl9Dnoq
LynNiHwJ6F2LA2EzrDS4jsiTgAf8MyKwbMTpx42lnIqx6IQiBf5+aLnff4gUesSb
yQph5F9Og6oPfJ80ths9cQ7y4/LIcudlN7F23aDbrzg62wMLaNTt8Bk92i+9eodP
9YP95UZa8Ww8MVPD8o0LfgHyG95ozBosTlg2Vxcw1jtGvuspXA5tTQu/l3QsHiTj
yUiuPSqgTj3gWM2VE21lehoWvhcACd4rDwhb5ckH5VUlxvZPiVONgvHW7GiVIKiL
fOGXc09WfVFFbfnysRr6y2jVca9Kd30CLtdXmCaoXghIq7IX0KQPf6bAbzeFbyn3
tBoAPStON+qAIf36Sn4s96C7/DgR/kpDSUp4kcYeUs6p2XHD0wN+hdgTRFOlgRnU
BAgGe0tIiEBKmCm+D1YmYiuuALvx86BrRFSKIr8m8nD1SXlyq0WiwbGUbKxb07gn
InPRmyHffCIQUNcPk13LvKJW2MUZqVeJsXRH8VM86Fu9FXEdS3eVBeSbBtmVU16+
RrAEQ4Ys9W9+77cwaCiwtJI43cC9kBj9ZDcy3H8jmwvGIsJ/XDENJ5Mr/qMUoWFv
+8rF3QutoaSbVbinYtQdwK44C+UWmqKJYQ4TMZi+j4hsRxXbD/+azjeGPI8PxsUM
6FJPV8kPiDMaZfEo+MGHIgrjsBio3Rhf6ylEP4k0NRDSueari93MApEgkI9u1ZnM
dPffewXgUKnv9eL95Lr0wC5rovPleL/28DidbVzs0dsL9Ybp2wDuqeYveVsWoJfS
OYFeLO3ONudB3GIWPco3hHZIv8ZtsCYbRW5+HeIwpuS9w+7kkMfgWzK6S2j52kBS
bZOPtAmfj0uX4Q8jxM9Yu1x5jkU/KBEE1xp+Xn8UJv6Wsii6xPRai8GneA6tipZb
KjVRErFRWtmHqlBVpRpf+6eds0ZDh78F5s5/gBG3qPLjsFju/55oqHYy/Igl3AxM
CxDuaDzPX/xe9/nGHptzU3AC1vUVuqxj/oSjcNbUw8/Hj+0urMoHokYllTGhNqby
DpSrLFx71cAXkxvN/5bkfhrrqKJwVSGJDjXxvf661wTMLth6fg2fXQqvQux3wlG4
mfrDdL0s1o22EaPGpIjIB56RlARz1dmiubopmpw4h4T2M4ORlXkecw0t7lAda/DV
edn6FXcxlZzxMOgmhx5LwoRQq6/U6i2QqxrvLh/nlwxWxDK0u5NFP3CqnuZ9lq0u
qq+RyPLjmDCkHHE27z+8nq2AexeTmXSJQszCQI8kj8lm0Fcb8w134LcGi/ebSXeZ
TIcWUfbBqOINuXnSfkTl8RItWNcNw7U3tVQkvGltYmvKhEXPkkMsSjRmXUQI+rab
u8d3gu4ewlRkLITUufMbRDWGfyegcyqDReDLQoZJyKv20jMbisA5wd+vkhlqcelW
73N8EfDvnVlP7alIad2BUD1VnfsIh0FuvHJgX4u0qmEQsWjh/xclP+GNEYHJst68
MhD8vQVtvJ4nGefIfTV6whKVsG5ow9qAp/40Yh64ZdQSgQS14jia3sf0jtFFL3F6
/1G89AGZ/Rxn+E6kMSZ6Ev7AGcwRzgWFEtzmkNEcgX1DLKaqwgehkH3xx17DOniV
8i6O2mj+VrmE9F04vhneWtOkKW1rzvm+eJVWeUOpjyZuVegg2T4nVr1oAfEXh3Lp
oCY2AqzcFYR2/Ws23zhaT5kajfnyjApNH+X/Uhmj5xe3EeHoqjmBu9b4uRIfO83n
90flbCSW4X7nQXJqFFv5KlTrIg8g0VITTmWifeqkg5Zk50HOKTKifngJOPWHsfNQ
FKZoFTT2HyWwtKwb2qo3M4wYhhiuC54oWTbTCpi4+4y05m4UnngCh4oKqDK1Keb/
NushGbjaVQNZgX91DF6g4Quyo1QiND62vPob7/lcxtxEnMaVV+7rzMLKzGG8YTlU
wOSpK3L3SbcQxj89rS8vHEZREhKxtJ/nUF9JxtsbiUG0CfS2vZ99pRx7mpvhcBN8
h/QBCi3u/rQ5hQleSpzZXF3evQcAHICfU2lbH3bPntupDPScBvObgg+CQ3qZZS1h
6/jBQ/Z42zecpmSH+ZPgSVJRCsOM7gyIww4jU5vcvn+QQRqr/uFxIcqhpGpcIMpR
/2gbQyTIQgNHCtmfkSqvysq2dr/saq3pQwFsL1W1zkxaWJacO6kXOojYiJ8slTRJ
4+tFAIvERB0sVBYfDyoHduz8TPsCsw+MHzEL0VmEJd/JhH/biHHTzSwrZSSubNSm
oCv/TDPj1Gxl50e9LD6OAlBYlUNbZORz6xPS4E8fxBsVdZc0BSJAK7tMLBlwYEj+
tN/DeL8Ojow4lKesS35iITlLfiBmmc3NS/hQFFYRTkFslMeAmfYhMoF8/afydD6F
wJRqsW3ndgIh9E8baJXi+AheClpN44xvU1Qz/G6+e/GT4FSlyDEFnbvFywJs0L7Y
78zI1dsQMazViXNSMrKhrdyy1rdomw2PWleIYUb2QXnLYFQhYbMvRr6zh8xXReTi
hVqzKSBmoVqDVpP56ol+raSrpaSq6VkJ7jBHza3iRgu58gUbUTJ8yangLFFkXhCd
WzsBhsuPS+vfLW9/zlPQyMuUfIJaF555rEE7LJRvMxqVMN3GlWSq5LbNZScM66XS
MGGAaiyLl10L9hX5Hmd/Gp8+kAydIUkkaFKaRMIlOO5N+MWEYVvdFBByRc/pZo/S
fW1f1z1O8W9SwtE7JBRagWZquwK8d1/4g5C/4MOvPdJGFvWDKRM0tivWwc0ITA45
jaEpF2kMff2ba4co4s448Yo1jcDms6qUMa4v4t7lOh4wapwGnF48VN521vIbY11x
Eq45J0Q12/OVxp+JCAHJYM+BY21CjnSNkzNSLBuv2UvqfssYpO50VjivEmqGSfHy
m7KFYY5i1/Nu6HKiJ2vhDvDFkrFoW076k2sTsJkN786GPtRNUk40nyrqez32DzRC
/W2wjqLM9+LF64t1W2ckmrZoZsV6NVaoBMghnKbgb8CRAkibGK08bZyhN+BBJg4n
0CzWFxvx/R6EEExtYcfoljSMo7IgFBWRMzaPncjFJLLHeZpz3OjJ1+LW7tqkBD/0
QopKZti43AufHQLZa4JF5zkgh/vzGJRSGP9wrjpbRj8MirRWbtiE8ZsTV4HkCYHI
QwrOqKkuq3dF4VR/GoN15PkySrTieHZ7ah0IA1lFNwYi7RGaPPli2SPorPa4icDR
IK/366xJOcTGLCOHJLPZvhnVj8kUXVt8nvVqJYoZ4gZz4GQ8P03OzxCcQ1NL9IEu
jixePeZ4zdVJUkMcgJjmAqgK2JSJo1xlB+CdPLzt7yauLYPbUdRSV3PHb0vPTTUD
hLnLE+8fJPiM/jzWhNM8DN4/5NDOvFVkFjF/EQ8y06L8dDnqLocwxWSSgsY59dfU
GZwFdoV55y0Y9zguNvFzzwPFaR7m7ymcjk49qd2nxMucZLWiC2AhLuRHPdiMxdcT
Cn2DwVIAIBhP3GtzY/V/depcsumvuP1PObakmubSvSOzt1BGwqz7lzDge+K48SJ+
RvsjSgoJ0Wk8+V72NaMRkWt+hZyS212CY8NW1a67M7gMxxBxwLqaPNpG9yX8bpXk
LdMuzefVKy1yJgs2AJpNM4soQqRdiOqjghmlanfm+5ccfOvq4VQy7oaLIhOhzJoV
4+EHuRw9moxs069+c5+o33JLgJk3fKIWV6PlW1cvQYGb6a00MYtb4m8nwEOmMZYf
oKM/wvckx0jcTNQ8L3dBR3tnfZGJDiD3u2/WNDnrZfbZleGxPHGUXrYvtRNIF1FJ
OuqDw9P2uSA9ykvLZnl+mZ+4c2/ud+l4f2X1kKokrWpVdXlBp1xIJl+75lw86nac
oZG9YSAtWL1xuoLcxu50hZaw23Rm7tOQuecKItBdqD+Zr4E7bKSVP0bphZFwGSrU
KDmc7c/M9mFs33QR3oTfhxK9iR7HxGHPJwbyna7kpNil190m+GYQdCbQOsv6evOE
xP+A3BWqsZdwH3mLct8X0g8hmp1/XPdpWWMLkgBRsbjOWGAWka4tLmeIZVz3Sk/U
/OQEJUdfTt45COOZfVXPmCH8ur1P1GfZsFNvNUYKvBPShC8UzZMngrDiQqupqxAa
MYgO/Cko2rwynISei0kZK1Y4wf0c+U00mMVqUSssm/85JMuFL7e53U9fFcKVHRxT
uZ4yOVHSweueDGJqm3AW/MItHatpzNCbdeFTaQcdXR3Kbh5OCG0ht1A1DM84H4bO
j5CEG22j2HnekL2MNiODdU8ZVnK1c9HAp1ncdTeX7zTYhJmIFSgpN63GHC6M1SGj
Lw4i62X8YTAfzr87yT9KFEUWN715hkL0CoESCpPjGfilOeXLxO82JY3Hq3Lf38Sx
y6MitF9Sp9YV+f0siiF/Ooj6LeujIOhGalRvCi6UreF1GrO7Lww3a5EAaZg9W2ua
rvYxhSeUZn0dEEBTFeyyfdujQ1ezbaopBZfgAwhKVgWl9sYD3QG+q/bFdhwA+hNl
V7RTxgZN2OchXyAXXItT3SEIyqgiW76gm2e2YjEbW99sRzCi2uk5hJZXlcXJylh2
fwpELqDMiA6/rDhWxkDaHaaPDEcOsDHg2SxtYe+gR48ZYcFI7eF82aMcfKcAntb+
I2C80frUTmNsQoO42ry+JueAyWmevj2+HaEO1oR88eTjTiPYbBsuZyfY58ypbwna
25QDNRvL5Wp334nSO3JKSKglF+J0Wd/1FS22/lWW5xHIOaEg3TxHsDdDFhFNra9s
IDuDCFExf1YJVDj4QCjVvPlMawzNQ9qdkf5XVD0B40RcL6TFXgE6CHesGfwI67lh
5l6YVQbCJGNx7Tpfx05VF6pYz598T43YZzNhafNoiwYkfbylaNe29wviWfXLGDO2
kc1f886e/PFQisH2np7Vi4DYa9uv81VL/gwL36VNbrJqd+YA6ddewQtXn/UFxpyp
hTtSvEB0oKzgZI0FmkmqUdmOdkcHXQhfhctOuVtcVbds5fDDNjv+btQZSEbC4SSI
GC2mdXCOVQZMO3lv/KyIfLlZSn5qEsYg6JMivr7NHuriSopDLXdYM7/8W96JxcEL
dVapRZAU6nPGI/IGTZerUV0iBQW07FyvnJZLq+hkHx/CxnxXyxtJTgtCXXseCvvt
kacj4KT+fUbX2e/m8j9GSREVKdV3BFYnpiWCGwQ1Lfta/XDMUD5UY89l/wuGSCtt
qKFCc8CeNvo8psg2itzgsYdmnYm99YxVzGglUUZ0XySQVTeio7Iu9Rz0vZo5byBB
AHsCXz/MOv23n+8idsJs4AG6syjvvABbVL4c4ChKninDEtvCbj49uFlwk+FSKk/u
dxcRETGMTytdv9c1bD0IvBu9ct1TgkzXDA293mD8DL8z12RXxHGvMNKk2Kvk9e05
fiTIZSP6dDjGaEt/inYpqlqNJv5QCbOCD6MdFGKGx33NC8wxeWLkA6zIsx0tWIYt
vhnZ6kvEf8sJTot4iBoNDmNrCAPA+bGkdzcst7zPfDZbml2o9bVTx34A5jX7XT0v
NcxSwNC1zhRO3pZh+Ovp7lTavaHkMuf+2zLrSrV28HVnRaSmUfzYPPHsGV/EmPXQ
MmUlyCi+BhdmJx++k3pFqDCoWtVjAZNjemMJVKXWQyKhHK8OA3A4XZ1tNbCFGrE8
TacSLlV83DoccEi36j1aWuukAt+VlIud9SgkgQasz2GEY7fAG5+iAivUCPzoWpl2
yWdcZsY6oAJktHEipaxsFSWLN5GpiJnujJ7waxwIJSWzpy6ByJNcAdmkAmr5lDTi
Vztb0YFnKojzEvmlPPyuDFPDuOrIRHSe0Jbx+K+hcMIur9EXBPWb7mfIoxLqJqNA
yQsnShSjL01bOpMWG4AxnNXE6fVeG6iifHPgEvQOkkf10oO3snT86mshbF+7dHSm
frapcao1jRSOgkVoI5f1fTFQoYsgScNkWu7WL7Ow5F/+H+nLBwMTYpoNq8hl/qzW
f+qNfx9xTDiKGF/oUEyVTuBIDZQjoPbxBYCG7FZAjKxD94APzDHe8uigc4xEQpaI
svbGVzZbOcfJpEmu8ANkc/Ke24XPKOy853RIX5LzryM/LS3ex1tQSg2qPjKDcy8X
Y4T2o7CwCVWd0ctBJCBJzk0GXuO6+Kx8KWP2deAmeeg5S0L5G9CMEvG7huEXH66J
BKNvzTf7m/uBdcVSnbvC4U224YKI9YCJc0L0lLn/YidjBwfWJ57PIhJO5bg/1UY7
Z4fELNXLWF/DRiGVRnillVkukAi4rbuVts/Fcmkw7CvwJicYuQQUvr1FXtfT01bZ
i7mrVK4wmR0heBh5wkpqruNS5U8N7xxljPoaq9+0eBU/BeBiiwcHmD4TH7dwiFWJ
6fGjrumto8R6u/iaw2Vza7zpj6pLVkt0YIPryXJ96JmGQOm/XP3DLuzMPRvoAHW0
kzVgIySYOTvUoX0ROXPZNTladTcJVVjJKRR/qzTdy2mXpTXCyrfrX+TvGXF1cN6r
RLvrzb5zT7l7vujl6mSZj95TKqdSm3iyJSNpj0i86Xo/bbp2YRt/aW8BSFDV53nF
JH/TzF4tTWOD9rEGExO9lhjGccHA3kl7jxe+ia+CfT8l+6eXeQxhyfE6bnlwSyeE
XQkiK7u90ZP23eisEC+lPz9qaIn+c0sjpIu9DWcsQr371OxnnhbdJRXoDdY4EpE9
z/WBBtTj6k8RnmdobYWx6GqNLK9wSum3Rc17S90uulRrqq2ojcdDAY8TtnVs6pZs
o4DxgLPHwK5SHk7WT2v3ZOCCfFQ8Cm2sslDCzrciGemem3JwrCGs82RusZXTia7N
SfNGT1v60rHtV5kLRJ8OqNm9L6Oc6qXWW6U6UOAkVbYj05yj9hXmf1oC/2/Aq1/R
BlAHoYC3Way47XizIOXyf1yGp8PbzZVwqGkT7IFWAi4/frYSw3NkTEPUIEt8lA26
qxo0m3vfeAZKLObaoLpU9nZLb2whrwLHsp8M1mEfFGkruZjBS5lNPryvnX3ImxeQ
R9kpfDiTcqYfnJEo5DCSe/+WkjsG40wf8/E36ZsKw6s7K1d2THW6DsgqUM1RhUOx
XofR+oY+8+ew0osdDByteFowQaI1PEVtZ3rH3Tu+zewGS7GP3DABHEUSJiaoG62S
OTZkMDk+jzDdkJMdAw5QEDD5xbRwnH78nt8uyPTyrQEWulpr1d2janYQZA9kJO5S
zZoe7ZZn8PLtvb6Qp9Qv/3mPAapFQDzuQ8BktWxk1KuHF8R6NO9ve1VCMvr2JIeP
2p+eZmP4Ouj1dtMITOV/jLBUw7IWpqp+RkySvVfKZlV+LtdMpL82dwvN4O1KnGtC
cJU6LkR1UNI0+hITEze71kJaA+R26KGwl47mYiohGHSWNEQYWdmpogTrrCClmidp
CoBZi4lNecAahylx0rxBwx2fR65OTiSBUh5XLWMRYfSAf+kJVtx+iXNdhq41+udJ
wM7dctqfIDgJ8gpxfbXT+vxad/8ZdA+5cscuS1BHGQpSqDfjCD3Z6elIGs2qQeJp
a3ee46LzO7FvGCURn5TBTAANvdmoBn8Adg8h85ieZ4U/moK8/k+GnCh4Yg9oBmZw
5iHWVmxhRbHGYfLPVYVEAwJva0XgBmiRqBzWO6AifqhFyze/b++gIhko5rJbAvbv
/NtPMDVaLU40UisHrIosqLFVu/2GCi4GsQIptwCcG32RJjX01rFs6svqSKH2QuU7
yzXsR/5qAVyPhfmgLuFUVqMY+jo5FtDv9R4tP9EUpyAQYKympg6GWOML4FsTGkLa
avh18chvdXftOAUh54AUYeN6dgeisC39ClhMqpIt2DC43LQ+bvl5cempzyWcIGF+
cceRylJmSaipEQvh/UyldCEuWweJgaxQwYWdpfZ/RDLpc+T5fZgB97Yq+6yEkFX0
h4ZCAdmN4ebhxLTzhz3gITx9bu7CwYHHM9lNgXKHQdrw6tEaZhvXFT8hYWVnq4r+
ZjnYQpyCpzgUttebNpR5mXHW3BlOpyQBFrY4uPu9cOamjeyC+WFV4V6P6W8XMAYD
UmpyjToR6Gi2xScx5MvigZuwGby2Pr8sVTdWy/yuH8sE3ujjULndtGUJHMDdI8d9
MW+EsAsPLQ/wdn4/ao1f2bxlnaC3rQypvTN/REolIIEegWzila3egBJ0tTsK68UB
aeIWkogRMZQE+h4hssSX5OYQ6G4WSOvBj+Z7hldsQEGMPMudCHb+81G68Emd5lBp
lLPRhWLAppRc+zcfCLZ/jVlqn55Z8fLfe2wGkUR3nUXFqgN3rDCPwTKafHY2EEQ3
hxpAyYBS2GdBOWSA4vC1Mf8qmPEOuFvQLDdZQ7XZdVH8MTBFnLsKU40MmhvOY8vY
yNNu/syzlUExJ+UnFRPPQvfL0jILaWd7PRympYcv6vF5BWHY8/hjg+ojE66a0r87
wYkocHv7ebF54078LADIOAbu7mKXH4HJkOWhdjS0ud9Ylb4TU7pjev8eaYbh5aHo
4pRYSmNM7+uzViA0djX2MX9NnLRuyCkUlSKEz8GTmQiX2IgcQoxP12pn67YKeLVc
9+MqTuxx5b6jgOs0MHNnCc6mQkN3SLGE4OZ59mPspGm3vk1R3JPfO5LHdiIw6J/F
anAmQZhIAEISoInvKWBie8fivDxNj8ozt5nGMVDOha8D4snsVCuKmf6CJXSBF+RO
+NrZ4+xZZ7xP5uEmMY0NiaVWkkVMyYFHW4rYTRei4e98KI/MONnPta+yJeBeR9MJ
/pEAx9aKSVfBHHmdO8uJzpUBKb1i/sok3LNruVom/3xBSmXtTKtjkjPvdVJ6QSXa
XSXyf0arglzkBCCdbXBPWBZgWvtJx68mQgSRJb2eak6DXqUkVk5BsLfzJCAhjN6Y
LbzDUmWkqq1N97j9dzrvoNqzzgOeX1utgfIxvmfa2eh9WmUBzszI3HdUIv/gb76n
ofPgq2o8VOxYoouzfCgNif0tpz3RyFvhhXv5HrFBcOInv+/SFQvDrpbSkfOSgosV
pvDqDLguTfbFf1DiJyY+Py+w9JsIXWsairVJkIGyWLhBvDx7eUqMJTHUu9KPghan
nbqpAJcnzWGZ0pcAsqehGEiLP0Ra7Z3yXbmEEh1r4RyLYkQ9n1eJ3rXknTBCz3dz
sXBovifoJ+Kn1xfg9+Zi6kDBooGyHywLB5NJCUgX+/QmxO3woaxgKq8AWGZkfT90
MPd3ZY400fagUofND+1Op0hkV6dei+OUHdJK+KFKOpSKbz6nIWpISco3K979de8n
aCzzGRQg8JQo+mlOySfGfITy3d9KnoYemBfOVfDU+hsRtI9qUT8bDugFvaqdFG8m
UvSOqTkoxuTrIzF0/uF/GckPZ6vF9U93XNvKSpgGnKy99MgUDueZO1kSWyZEzq71
GKe5N5scnx2jf4Ym0N6jIKnyONeqg55bRbnqFE6d9bC1XXEgkinf4R+OkEvDuf52
WB6CS1uPRmKjmMdsIcusY2Zzn2zzXuP8MY1ktDLG62Ewvhst4m7/y89i78voMzkM
X5rnJYO6xSnh8S8DjmkX0BvYJe7N/OWBBZOtmeGwCrms25trbuT8egaaeM0Vy2nZ
JXnASPKlmCj0Ml522BSC9MHYj9ZV3ibgTmP69QM9FiDmx9DoxgwPRswA/L4lUpDZ
SxSogru1QTXG5UC/UsIhp4v5IoKBdQLSv+3qWa8J4MfDmawZKDY2YvNK+m+P3FOa
fuZ5aATLL0XbKAhXg6ZZBFLRu9m/t0PNI1Q8q9UHdPKJHjlMWpERk6cV8DfqlW05
6K/FOfnUjifht9tRRWn6G8t7TDg00e0oEG+bTu+BVpOybql6Xw8yKjgHta8cwbDh
aQ1/DClknMQsVxghqQb4ObPz6mYuLln6gDJPTsXXMkQUc/wObGf6ydh8v+dgU5It
yXc0Uql2P1SarJBEHab2bnOnj8kYyBqzKhlTs3PHtdDB6TPuEytwSutgN0sf94k8
tHYKS9MOXUg/BVO6C23MbpjX/TyrXpqGh7nMIulSntfygpa6oVCmXwmkvUVrlEFZ
i4h7joUhGEBfZapOipqPHS64DOQEcLh/3doaury9rvZj6FhtP4k0K1yv0cMPh4QD
DYTZFoWI2rms1d4dwjX7r0H3j+v8znQLytFu+tOYUXe/PDOlAS7bl59p8pVkkfiN
FcmOkCZIt40hx3haH+h4gq8+O04QymFDmEREnOPNYb/LcB32SxYb4NIwzaO+zeQi
jY389nufqcB3jX7/vRowgS68EaKm4b2EYuT5MI9RDJwvLvoLWKZbuU8ETrJJEDZN
dPyDcA+aebCtMp3slszIMcceJdRcs9VzSenn4gO6kh2hXzk1SNYh5ifvkjUnIGuj
XZcRH4JzPNL68I4dB5Ty+phFJOBADgrX0C/o5212AkTjPIRvkaWnSFr8z/jayY3g
N83M6kXGz1YZDClwreLr9g+3aInL0SF2Ffmg4eR+1+wFfYjIuaiRemBjLyAxBcSm
ZFvKTZwXwxConEMVGc/CXDL9GYYUPpZrdJxoyfYqLPziu4Z9NnJy7dU8nZ4YwNNL
kMvewb+4ipXZETlwWwd+uMItJTijk/++ulHJGAdbk2lb5opnSE88tgsn7xep/05S
Xm2S79tzozz4/RYdIt6z6yC/RXXuWqN8QyQ/ozG3of4dFHWEs5ToK7NflQEVW1eW
KIm5UhnAQf9+YHQgNsPbuZUmDSJqg7J3PtrzSrdUVIzK5BUxaR+GsIjNzSPea/H/
H2Lu0ajp2QGBFfrzHchCFAYbE38JxCYGzhWYuy7yRwnSeVTM7Atw+VBaxkEHYVJ7
domXJdKdbRgL9sCfAaXmBZBHbO1Iz4RC1Gif41jQPAbRwlc9utpAGiSYQdmTdJkQ
EvYAzxh2XWl6uIwGBvzH4FleHowdlroFGdN23L0DghcIbkzh+5HSkW/CeCWIjqFb
7PbMFLT1xWiLj/ewovoxUtjUs6mw4zRTIlvajmm2q3IRA3b55eZ2qCBbOgBklLup
4O8XNwBr59IvcNm0hp1HJ/WAHHdC7858qqsaWWWGetNzAD5QcjqYxsuVDqinL2gf
zXL/GIOFAwfgV6s7zP0SO2dTRHXM/VMHROUsr2Lmx9f05y93ctltMBz614zl6dTH
NHeJcs36wVexKXe6ztpTF7q5YhbA5687p74THNi2LUNlGHtJ8b1njvKM1L14o28z
Z68oF+izqub2GzOeQmhRNSpKaQyK5X0Fb55KSF3SO+lu5HM5VZdbDss5HF7kE/z+
xdW/6uMfxbCm8yEt3coC/VX+2S3ZhivDn4+7WrW4tcL1IY3fpOM+OorEKAYH5jyP
gSq2mezxv3pHSGOH4kQNxGJgyWJjzqRFB9SlrQUeHF7vIlZfn/xcQGZfaPTt12BV
l8okQGEu1j/sc3v2HRCmFk1VhjVPKpOqsLQARh2qDoKQayHjjKD0o+a0rWC0K7ka
zfNnb45vmsqyjvnGvqlSLxAH4XlgFtVN2mzs2NcRP1Y7G1o9p73Ysjrpa2O+Xdzy
2Z+8wdveFnreqkeFZ36t3Ul1t4RKWm8oJ9YUs/+bXcrynycNdGSnCFAa6mTpoukt
cm78HVPyanjiPTYES3GozcLDxSQIOtDSifLCNTOyDlC9jS/BnzHxJLfSl77Fde1l
d7l943hhNsUNbhVWywHcHb8FVXqhBRc54ak0EIAjaxB9KF5CY4LNUVtQ4eTGeT/c
MuSGAR8pNGA4wGDAeiaUEXzEh5Z0voWEEmWAKzZzqBGGce1NrpuOlsGOGcNXTCS2
QMzmIVsB032nyOTLuJ8m5akC+dhLDjYvXOELVdzGUEXeRnNlQyyummIRjWEXXnFL
CtG6HppQyqTAlgZzYwMhdSJRrTaGMBoZy0vwafXxbAj7GK6jijNZCSWz3t2Y9BcL
hMMSV5EEpOXbfRhsw05H9ZlKspXNtBchy16azuNpBoR6YNQtmPxnTuT63ubDglgV
zBDpgXEIo1tVM+B/dCnV4wZGq6/2Lc1pl2r32Qprh4ZKTQIoGSY1y9iAYisSaRRF
CIPtnyzB9grTYDlHesiAKT/b00oa/mp7lflYXlxqUmnBOuH2LDHb13o4BRG7epLV
8EDPm8p4opygG9g4lD9i5ppXEuW+4ENnpGxz5ymQZuI1G+P2gllfvfbN8/e7Mpcw
goBFpqV5mu8CEYOyVNPwRqvNas4CaZThtqD/bpZqqIbh3sGCb5IxBnKwQOXGr5/O
SSnbDMNxzNRqI8yyAzFV5os+6mru3jyzTKhepeKD9yIdEe6uGQiiZ+mpbQnEfQnP
LpSbbUzh5ILHV15bIwfgeWGshHwGYZaCMUEwYMn6FcW6Ej1zdujUBpS6YK1DCAgR
KQx3TbHlGwaY0rn+mzbzx1+3zAJFN7UUlfhTswvO7yToayb2FYLpBWqBg/4nHkPH
zZ0nP+QzdrcBgBseuPOk+tDwjW3pgN0ZcjRtFKwYyd8K5GUFIz52QsPdvzZLr7TS
zuLHer6FKt9wZpYotwVmAYgyFBPX60DvI6eictGqCRjN3lRf6wI1z7xIwyNce8y6
qiehBRGWD5WnK4BE2iVUu4/v8q624DDStSGTGp5cbh6ode+zEDwvfvFzAQi3nEUG
RhDo0YXGr1ccL8RMF0R9/vA8WGGn1mUqKwR+V4piNDcNfCXdvXco6SOKnTBdWdeV
1WyI2e+HgRGWNSecbalVuAJ89w8s/meqDpJ4gXlViP2++t5BOXGJqsMwHBgzN+o/
RF8fzb2cKChydhdzsFKBrd7PclK9n13j+r6ve2deFRfZAhk2cX+nRjEJtWRhNxVq
pfSDHvcXfyBWXe5SsFf7oLUrsVmiV6tzFav4Z23s6u1KTbfF0GXbc4Fz7J/4YEr3
q62VgWpDf8kxEqhxz4Lts3UIOBAmNf7y/gUty7D5NZC+GZQCfjSfkALfQb6ROjVW
j/XM2gHB7etV7eTIEg4PgcgP2OmnYheiRRT5AO29fWyKLdRwAhk2pwQFxYxlGplk
tKkiwEzHliNN+2UZOGaD5x9Xzdrgk2UKggsg38Dl9Cyf1dr4s1iA33J0uAdVuaTA
9Y27RFJCNfYkGElGvDMhuibbAgpsIuL8HZC33AEDVRcmCxAnmqGp/Exc9YuHE6xe
+R6pVbrru/6IKPTWJ/eCU+ev7HoEJzs4Mlsg/HMPVGnTWv1QotEgwSVcvIPCx6/S
634X+iR3vGIHWTKmU3UjXv2/hoaTqtGhNE8vrFAY8Ci/Rec8is6SAWNLy4dOJoFY
gSidbZfi3ysT2zjST5dVOuTiQDgZZcmXXqkTql0AGWXTzYbU2oYGMP5glaWJs3GY
s1MVRMmYoz575y0ZJLUzkeqOXPgHQH7gInVTKSToiY9vsbDJDxaLoXPm/QEOQWTR
zjLqe41m2VA9qfERRzm9cEmAgORqWI4ub1OjxWu3uaRIPdhSgxiXQnQSz45sG6vj
Ve/ERPM66kTdNseRKjC5nPy3fLFk+nfKNIiRh8Dl6OX57Icjnrvv5lGXEReNhnxj
yxeDAU2upz7GjPgZb3kyFzl8xdxfpD7cMz5FXIYHZmhDL4Xke+XTpWAnlMw3KbEL
sPmD+o8RsmL2mwgNOfP3rMOAuFnenAjagTzykWsBM1o80VkF/jKWayqJjsWRZSUD
kZNRZu6ZAsYebNsjBbo95/T5kzd3O7YY5GB53QLI8pa+qLL0CuaO6Xw2BCFKypzb
DLNvN2nVmlpq/xBr8+NFUMJ3myIZSNcayiunzxKTJsLxQTgX+aKZDfsCLG4cOHcX
shB2GNiDKCK2c1l0jIjk8awz6OBH3InILq6a8y9RmkKXs0SfBcYJxuP0q7u4S1bC
Jdj0iJz0jat35DcSANjv9P3ufjlBHrKbZH7TrTPhuIclk3Y1XNht21TyWbWAgXdZ
di82qLMv39pn/8lyGEt1Ba+H6NNiwarHoYTFYE13Ex6liEM+UhkNSY5fmAVywz/i
9KkpJBd0Q0RXa5/tzma+PgAWW8DBkaQVxdRc8MVea5Jioku2PYv9cYeKiH4JKnie
1JnNIVYLvdqq8DN4GurVZdG7n4aHvzbdpLMfrpCXPu+fm/93cP0I1CyNXba3TIXp
7oe6ZCwlhjsgvYB6ycwRS5QiZ9+EdzGDyqrtHqljMvsGeng1RrTeEhWhsm/VTt3e
D/3L20wRlD7echk5bdbgCY2xANEIbm9wuY08Oiw1q9Xbwbbaxo+M4u8qEwKENqqj
c9GlFmHn1s/5d3xYsFBihsdA2EqDGNIPWkN3r1mrm7qyH+oNiTXcxsLjSBoKIxEZ
QjcieR1oZdabeoHO0WHvM6cmh3qfgVWGEZ3/iE7HMFxicD4Kocnht7WnjYcaKjHT
EhozFh7SSe17ykPKVPFrUrhbZeG7A1b2Ys0x+GBGI6ijY8gN/Hfu/8CSIraMDdnZ
KYDrRbqzbIkA3v/31CUpaJmV0aPfoIyCDfkSYwDk9dzrIsFoUb3+BnaVT/l/H+tB
yQl7enPph0ey46YVlpOw6fhtmqLc0Nq0s8LCPnlK/GuCW0yN/GZUCkt0nCTx7V93
ozMWd9N4DZ2A04nDtDyKNLrB/cqCqzfFtAIm5G3bCGW5OC4qnI1y39UAVe+YkeAJ
emyXf6HuYyNZipqdBO5+8oQp9j/QWq2D7LBPOZxAeLXte/zE4/CUZ0iNGaBh3bvg
TU4bdrfIkULqlaq9kDJFWLkfeFGY3ynabgPxQ8HbRQAK3ZC0+vUaRGnZnSWqRuyV
U5mlOSjNN/1Y5gjcpvf/HWmoScXFdc47S7Ig/IXysjuU7v2KKx8L91RZE7zdOm32
qCyEIOd80B2aWmYuGv/e9WKWfWouZhu2/1gR2UcjCzYYuc1EnqlItj/Lp/swLf/J
5nU1p8+1t2+pCAcmCzdTVKYt9r+Da8EIhVdixxj2C/J+yGe+kzB2mqVKJ1nBH5Gb
oOlsh4zL4+AMHWfipc5bvYfabtJkd6mgmtc8JymHjTcVVDGWYuUpPEiDEWbgsEYf
8nTRbB8A7leNxjvf3EmokZD4lcEiG0dEcn8B7moyibafgmfYlz+/TckDlMbeme43
qzj08EhkSh6RmqzHD4rtoEA1fGxOgnCCYiTh0Weg43bpRLXIilAHAEB5tSN1Tn16
cLj/soeGCcdRX7BsD8l4HWilcFZXeMmZ77z2ElaQyqBBXZVEoTRNRTSnzkiIzzqk
73sCUAER/f/SaNPLScgYSpnTT8IBk1nVy5B3A90CHJeFixjANVzICm8kBbNbMN0m
lqGhyBfYakD2RSL58Ny2q1c3u52Di5aksuNsw5KLv3df7Rk93wqT3TP9GqVwCCHZ
Rwe85ses4A7Lj0ndKahqM2pRxFmRPbMXT4IqZSjSB6QN+F/M+HflaDihETCrW1qa
GkUQS7KF5JVlnBvwcFFUr2iOe4HhHkJsGbjWo1ImM5HAAl9q0Zqu9+E2xhL7Answ
HtApEIjL25ylRl1j43rWZETHPhesc3OZqrcmcif8XLBkGcWzQhhi86LrU0DNIIIr
oAVQDY+XE2cs1tRQDKpVmjuGvvAHrvzI/knmYOAD1eUVILfDTAuclh4Xw7DCaAkN
kMz8dETm6yTtAyYj2oaz3y2WdEt1cI/FgwuvnvbF+/XVj20nkx9EqUuH750nOKXk
wWqVx969Tf/H/CyhFjx47I9mbLlWG/9fO2R5HSg8mGasOZkr/fAWGn3d4p3CIP4a
oAXz1110+ooLgXLoFXo+FKGjqdTZlOd81TbF57MKDpIdgNYvRh2otZzI5OnERVgz
N+r/XH+5zIxu9uDmOdjWcKbnPn8ruG28wd4M6+uMUMPN7aTX6Y93VONOG0KDZedU
C1BaLzwbTIcTE/M1wyyKjN4O97wMYrIxeGxKm+6bWkY6WJoGZV7r8LNnEaT7t+Yi
bUjUBbolgunyAOfMqpX7yf7vZG8xdaMVJvsaWBemhEE8JXpOoxhNNy9laSbkpAVj
75Cj/3OK9k0MsqIwroVS9MNuZlfigejdUqqc3z5HFzuXTBa9oSJPWG6FKFhYFRlF
Mq1d2DyFdTt8WDRYJvFB2yJFm7MV25XX8QLbCONq1mGS3A/c3X1clq2ng3Q6c1Es
ES4MMw2/FPSJeB5U/I1OyrrKowMIWlSk3AduYch96PuI45uO7fQXDglJ3rv07xJo
evCiMa2zKpn09goaDozB3E4j0OwxtRAirWmvd324wl8N1b4cYbZJwKJVpRw+RO5x
oowbfyAagOqR1nbKxYpA3s5dnEBTNeFEVCP21/xHc83yNNAk7l0bRAWcDEKaqezN
QTYiKu6F0Bxi0kBAYwd6bDTLW2fRA6gN8PxEffI1AWgDGFfL0LYVKG4jhFjsnhE8
iuehse5KSG/6WlHVSKq26PhSVsh+cMl3MHH7zluQMuryTft5/MVv6L6ZW7OdbrGu
YL62eKcvu6iCGOqIHY1KmsnX5oC5+Qz6RTyRrvaQru9U+hbzgDEgw+M409AjjLmo
IKEjTaCVNPwdrK+f8UR8jM9hsvu1yPu6ljHt24MZUBTWEn5vNu6VBlF5RMB5nE5d
6Nc6dp0MJXvHxzjIUaXyDRwkwWwxPhIHcDicnYNmL4T3jMviHw47O+gKL/kjSJKo
o8ci64IjNKk6JWguIZLH1sCa8haYkYbX7rRi6vhZZw+R8+Rz7cC20R7ZlkNvXOG3
nwCPlkCJWzEhLgCgPEdcsXZpNt7jWMCSaWs9NVTx1ALE3X90P/MMkvytqjnfi9Ew
w0+Lv9sXhY8FrXMiqXy/39h6Vr+52jpuEpv7wKiigMbtp78tgPDW25fAaF0S/hDs
NVJC4tq7gLZ5QNtmRqgXIt5Z4tCgIKsQApPdpW0XJHEKjV5SUfWTRkvb6fqdoupZ
By7olqMXzCkqoiIqEpm2IBcDfZQh+jejcZ8KNFhw30Kn5QbyPc3EVW+0G3hY4uFj
l798Gu0/GPgKBRhFpRU2+rhrv5OopndWlbCdRS7J5AnBT7UrtLQ5dKYOHxgtz1+s
cTH5Dul4iIbsMG9WUlfFAWwgVYE1HfHSU63zvlvuEpJcXzdivp7JCGr/W8Psm9Rz
xO7ydvYnKcJT2sv2wfMZskaevb1dO/bqIc75wtB86o6KCtuV/vtd82hv/U8B2X7E
caLykMr6Ihxt/3cG2nkWrKKi+dnVNUAzyIrXyrOi42JKn37PWEbfKkEiS/abQbdj
Qm67V/PeC6P2/Xmpx0SBI/Oi2YbLsJPBsidS4JGMsRqYhtjS++H+cFVi2XV0Qtn0
S0vMizCxwtI+GOGdfmMLKmrdRDo8BBnMpYsK00VCKU2Yv6ErM5eOuYN4q7IqI7K8
OvlVNGtpuzZo6tX49JKgSOU21C2HOQ/Xkpoq9yZTqYX9D1PnwE9hlTowQYMZTxjU
clvlnRUxwW/l/GmOM3dU4O5sxjWHYBaC1ODzBrM6ep27um9JBYAH5bqoCyiYEMa+
wW5P95CdtIQM58pmMJOY+BqmGblw115r9R0AvqcVEk1ZcqEX7LWwLFZE900upnQ5
IAc+du/pYvIVHu9PAW+D1d+VDr1RWCcOiDYD/6DkiTq0+HwXjPhvyibZtgMMZso1
B7JrkcqgAhCvfB5InAvqQqWBuXJPTv3DwaBaak3aPbw9ZYnROkE3l3UatTc3+H64
5jBd3GP8eQO4GAGdXADSV16SQNG5UKfCnhPngzoZ1fRIioBTPVvHssOW+aMLeM/N
wGXioJfItvEnpGrkfWWhO0TfmjXusfUlJDk1bffUU/y/zCYjmTeCHOmssJNrfIy+
JOQm4+m5Mqat5b3Vrg0Z7FxNlbmvGmfT1MbHaqNWzAVwRpvSacUIP3ofKG44aNq2
4LfEhZ+oI41KZWLTm/gKB55zkAEw/tghAFo5rNoo5fJvp2ML9NOGeSkPPBIVJuef
HegGqZ5UWb0aV9unsUJoE8AqEEo6Hoh316xXpn0qW64+OesqVHnGpJChVtWuIQ5c
E4aA6G000fI8R8baok0PhUIO6dCcm7mPdSVkZazF/sbxlIIPChfAug4s3mkG9HcC
0yVaEhu3+UdOuvxSJg4WMsG4ywb7ETlka/Iown+6pyujnQsOz0wkfSR6epXFB/g9
IYkkmmBqyREIsK1dXQ9M74VR2DAvONGz4fb2PknGj0unCm3BGHa3j+a/6mqv5mu6
TW5CwFl8rJStR+7q4bv8yzef+BSzvg0TXUEvy+5gbsqRNk8l4OOc9oekyz2nCdc7
M+cO0TsCj9xtZBy3111ECON4BGt9iAnYa0Vmm7LbSpsJGopfH1oO6kJeZJ1xRMzu
S5rlxcSbOGVlieMWUOLg+czvTq5IvvU8pyD8lbPKs61gCqDTd1I8nMm9j4N2yUK0
D8q1EKkjsTV2b3WMDNDPFhCbKniicvxNLN5rZ9S+YJnKaL7qwVuaf51EHjAtek2N
vCJn65NYnkdKhGKDfQd6Z4Trnq4ArB4J3IEgbYaqQVZy+p18GQf5P1ATmQDXKkwT
HNaVGOy0/INeMLip45CTXZJgwDXDUgVJCG2d9yguHfOQh2grziCVk0WorjvxTOtv
rVhqtG4sX9jzpZe/wtyrHypnUTe/0FDXvIHzJqFfeYh/pReKhtND//OQNkYIO6dv
5MglOFwUPjOrZZKlIW4JLHZqmkeF7a/cJWWbiyRr5ZNPcJkD/RJ0tOCoUSkr/6kX
VSzt0ncZJ4hlK0whx/7gv4S3PJTAevCqgcpKNga3SSbtWOx6c5r9zA0rYGGnd1n1
vFEkbBNO5/ZAiZ2gZlbO8fUUbebZUuyPhDNmXmQFFBosYxGKzCUpQTe45c8lKUFi
0KBPhbCbcoudGA2uISta6YLcTtzdOnA80NRRIY8URb2u6YbcJxdUnkzDUD14/YT6
uYyhkZLBVBPMp5Vyp6tbTZHJ5wdxzbk/+uFO7w4d/ckVcrrk25hRlFxRH2RZN3dq
Qt0eSOe2LZ3QG+xH9hI/MOAlfioLQa6AH6cDSoUlq9YczrYEBJ1a03NTmoWTVgWe
feJKa+oV5bgnyL2sHTXlrSR1p6+5rLaeJPn0wtcEX5tA3CNhdJ1lbZMv0uXnESSH
EnpTCgAXzl2/y7+ItN/vc51LJSUG9acVEzXjowabl16WHDHo6pQpnFzOq3shcolM
1bgxndz/WWgp6dwEfrPhPYGRDmlYAoRlhKl6IZISJUUXPQSQVaSDs0EmLI2pBeOB
zhZ/Fi9XvYy6z302CGPHmjcc7lUF1gPxufy2eQJQBo5XabuFkkH3oAkfIcLl+I7V
KV3T4mJufjLGb35TLhX/WMy1z9UwEHWWQc5wlRvcWX024JTOWKK8XSRcBCWRBFkA
D1umx2rIUUUS13F26HKSJPC06zO5ha6nSMItAKXuBBYRO14NASBrecJS+nA37SwI
R/S3IkwUZ3CLEO2P+0nqjmO7LEg5J2ST9wXe7E55h57+1VIy2tQ3nAK37MEJgHiH
wZFjjQy3hN2kN7jx7EPOxdtOmWPrT8Bop7Q2MAhBzw2qZshcz7ebzAforIqsde3d
VqLSCRQYZcVhQHFCJri+fW3SIP36GquEQTnKz0PUHRf+TESuQ/M9Sv3ak/Nt4/VH
p1VNlaDpuXNFJZypOTpbCoSda8qNHyyAaABMb9j8iXVWtQpXLOj43jzNWSPv+c4M
q0UP1LnXpkoCpvzw75h9+kxsIRn0ViV6eapMJ4zev5yioLCWdBqt50vpwM1OqI3k
UkHsbPj410m0FO8rojV3RyFXzwOjneDqKcZX/H9idmQ6j6UEFk7MuBVzbTW5sPSq
SOGX5EreeLLqEaxT/KC6xaqHJlVpoNFRwtOfYWWfjuxtRuiEmXS5aoMLcVRHW2cj
2F59n4GOuwbs3Vgiyz+Xulf1AOCVpbrXW0kTLpX/UOJCpLSOUnP83UnfEgLQEweJ
dHk11Zi7Iy8E7Ujc8/1P8VGZXCv0e1XqJ0Ss8w2TqFzqQSmDjHrYuaAX63jUHOXt
x/uTQfqZMfzapv59gTkA8OLSDynynm7LkPfNYdBD9UhQ+d53KEpXYfOmBJguJ0hG
92JBiNWePp08+v2ouFtIRyRtrWcQrHJzgJknoUk/pBAApwywktFkoZfI5SYoH2V7
GwUuu7ezPyKnHTbv2Qm4Cd+y9N1DMkltd2TmQLdGXkghL4MvlBnbfQUFlf8KuhLu
FL/nv8PqsH22fjBouo5zRuUdM5Pi7njoa2eTOLRr6LLXm+d9mpjRrE8RjlBtlZRJ
EPeU2q7s0aiE5WOfenBVG+scQFwOOZwNDhEUtXGYheeiES/1rmHrmc497KlGXX/n
WYmZBM/HKQwzqN3Yzv2/Q9aEmzzyUzI3m5P2bnK1+lnT2/YCzb3ep3rlMyIDi/YT
EFDZj3FqcbE7FDXT5gX3ped8Pd9YPKoqduHgNd74cQPSCasEPvSBkVh030yrDgF1
8IvluFePFSmHiQmT2CeazR4DSImkrDe6Etgo0ypLVTghHaOdsyM/L7xO3nPzWIwR
DsOlXcNNn9FQ+U8OkI5WRDfcEuB7EwOT3xXIuX/kut6kMO1dwwcAHMS+ZFXBKwrN
rz1UQCTKIQNVjutJzfkKWOq9Ew5GccwxnrP8fnOO22VO8NkWL8ceKRgcnxwI0P/3
tdOc0BBfRi7z5IG4OmbCA0JeMTOUzkgE6pX3CuZv2Q0INKrSJb7l4wB3EfGzfbUm
PTKF2/JIVt3zaOyrBqvTuk/E8mV2RFyU1mieXJmmSh/4goQhAuLG9UykwdPwNFSv
Un2/fcysyAWVaOFGJupytEdv5qLWbV2h036VuLKhpADrskwZyqK2ZfpatlqhvhPF
Ka9hYb+XagaxCNGYO173TPQKRsLzofX24VZOx3dtqZ0yXByV4RPeYmgq/9khRaIk
XLZjuhyXasq8TwxqoPGDeB4xs1ZCYPfPSX8fnrt47h1rd+Xtq8gFURas+ehxh0KO
4+hxgYThLUTaMOcGmZHGWaBKo2N79aPdVy8qoycRbG6fkxs1PxwN97O8G4zoPYw4
Jci+u6m/m0FUfRV3db9zL0zfsf955w202cq/qOEnBzgdC9V2tfEmoNei6IwjknnX
z82NxIKJ7hlpkL4uDUY++8k8GDI2kh7uQYhLaP3+10EkvnHMbM4XG7uDnw1pJ1iv
jDxDbRFnInrYx8+ZMeO4/Yj7Nt3XTeXj3qyzxbcszHD8d0a9hG7Y3Ad+8uBGrG0c
oQuENRNmNqzPhNfv1UYT/ncWofASa69VpxN7O4oDB42NJ3Ggk/ne1ePtN4TCiARs
c9qOdVcAjfUnsP9s6rDThZ9RhpwHvmXx2tg4GUBiwtjyo/dFO6nvWpEdFiGUjz2K
CJ5QV+Bc1RVSKegdpCcbblFbstc+Z2DIHz5UPK8R/PG7Ml1huLsuj7umm6I7UfpF
+zIwkeSdbQDrk058VBEthN14wifwmSzGE1hygNXfF2HJbJ08flPFMpACeK6njT/z
KPTU2lTdymt1RvlOJ7el2QFpJBPL97mgiRwlVbExOYOYNegTci/8ruHH8oziYKd9
kAdxWl61GkCdSyMLOBL0ogZF9GjOFdMlTaUYKFimeBS6tK/WpQF7eRVzLbYaIqxq
AP6HJEXwcVMNh6Eb/deawpM5KnE9b9pbSENtoJH6ktNHc6UmoEzzz6HAfzDTSvI8
FUK2J2iVpAAsxBgG0hH74fxnYTjFqFJo+Z9TjfYblHxJ7qb6lERlufTaPFhi1nQZ
PTN06dmEjm7mRuSoZf7x8LIWjaG6bT0za4ZmHusYz8ah7DtCrGGlPm9MIp/WAMXL
Gw4obaxXk+r+NVTZb5Ws34VytcBEtlwK5Qi9wF3d+7w88RtbjXDLqu9zg7x65hbC
FJjjsXYrClNunhqABgyLkvVQnQVetYusnSTetxmN4heKf+ZtrFRFcs2EvldQog8W
NN1u4fww53btnlAIoH0BUY1fKCcl7wF2IbBoipJMXO0k1gIiJiQvm0COI1H3S/jQ
YNFMTyPWwD0FqRJdNHhuvDfwksXK1YaFTpRYaGyJLXgiGoxqpnkuJoGX6MKP/UZZ
Ip89V1yhgbKJylku2wcuMFFM0JZ4tb+TNC1jlU9IKT1uDUQTvXXhfDb0LTvI4w+H
YAzBO09RXujKAzWQPqZTUVtBNamDSPt4Ttv52/1NF2+8xoM2GSzokPFmkhr32N7C
1+dlTTzSoClxy20RQGDoaKEaa+QqSNgXA9D3vf6LfwM8XxTV1+LuvfJfkv1PIRdd
2Jchz/WdMkXPRyhC3dLrhF5YoyeN7Lh1owV3nipuYxp8nvkef+nL9/T54XS1TYnt
kPgi81SLL2Pb59ZddKBlnlivC9zdtgh1kUKa61UlrziHVM74ZMGHbUAtLypd9SwA
GJbc0+rIPhXzMXBlG0+XuQ/uC2vYtcH1DAGgdZ0WI2yjg6MSDScYDt2hEapI7O5J
8Rclk9mUFhkJGVRDctT7JiztAMY0S9P7PpcY5TI6ift0YC2wn2v0JPAGZM3fftAa
d6sAljzAFz/9kOiBE4gCjDgw6+XXCzQdFiJsVBxVZhaoH/+7rOvX+JDsLUELWkhD
v2+2bOYGpSb0LpUGFHQCqKhpSKx3WYHJkeW448+yve4aeO8h6Fp5KvtBNMW2a0YO
J/K6A59g5lEUFpSRH2A/IwNtz+2NHyRFB2jUossQKoJe+C+9MgDqyK2M6kN7XkZ9
1aB0XUSPCgyOr3TcrNJG15j7JSPh/T+2BAN4Z7DEFBm1hK/y8C1IfNiPLa5vLMtk
ABNb7PKnqHgyS7dhiXvnCbMvHfQNjVgp5Qycblw4IOYLV7e20DpBU/LpIJ7wNdz/
/wRWKfVjjJVXDganxIdOV/o/fOElGoqEl5myP1YSWqWFzOm1jnm7a+Mpxp5KdvuL
WihW8Msk7iebIw8AXFbt4D5B/jGkG2IFhcjebM/mCypLRnmqLOzmaDbGxOLfgFZ5
4iUWoItCrDXpM3XpNsdgHl8szr8l2HmmELeQVQ234NASpS+cz0tJAAXKYm/axvHp
3ut78Vz9ho8Sgka6SCNRDdy2j1kfGWawmY2YjFaIcLpx4IvgDjrU0S3iwdpRsyzx
2YoCmjK/W1+FxH1WAItSNoYkhswPPRF1pMjBI6tByT0VsA2gqB8jRWgo9Bw9Q970
VIiTQGWyNJAu9NAGMIpQ+n/C5nyoqgMsYBYAS6e00i0VBqacN0GC4G5/RQmirnkf
NiZ42BzZESFU6Elv6Qkl48eV67ftNFuhnxMRRrguKgPw6HotmUdu9tq0Un+XakDI
Dh4QU09UvzwcFSDRa5Xq5oFFxMU/muXx3WIRIoQL6syx+ZzPD84SPZsZhCbEWcaf
KA1+ZNbmmxXruIhkLUcbAHtTupRdjDLAsZ7CVp6rNAT1xTdrXTqWQs4uFF6FONh3
Z0gTYtgcumfDFtIYLv41K74B3aAuyqGgw8N0BTiaKoC4N/7u5XEWH/4jbpGMg0SB
o0tZCjS+X61RZfiBQLjLOLSrSlHY4usNE4jw8Yr+VW+TeV+HGfb96CwXTWOK0MPe
JvCDCWY5V7nF3yfE97yHrjVHqcNzN3RBxr0UQyYADSFJGgx4Gg9foPdZ0MH8Pfl/
MAhKayavMfxUH5Qi5zkhGOWJkYTMJXhuwKMBbgfGs/iaogBDq9JWpSTeV78wsLbF
l/IiBSJg61vnJbxBJeWrji+FNcZrim5aAucVXXQao1gjAV9qrHiwhv1E4iJHVuj1
49dRg54u4lRCNYuuopmUyxnUfvJM0pTnOd/yqGVCydFhkO22Cp/83k7Zujp0Fz0X
qq0Re3U+10JtvpC5s8Q2M3nNmID2+kWMKmX3OBOry9Wp+yp38K8+0q92TRiCXmHv
DTv3pUptpi2JZDJjXlsYHJgxdPqexEBePWOxFAcwmFn8OTosMjKwrPsMH0zPcK4W
asyZEbgkDGilp2u2eC4/s/pklYLflzU5bXimF/tdef+ZkWrj6dgc4ykKWcFE4XbP
o1aS6hdijMB7wsfvnJj3zHN24ropOPVTWK4HXWnyb117ZgTj+fqFl2Rhbcxik4Rr
RxYVCH88OId/HsUAy+8t9GT3/MvAsGPlFlIG3NfbIIY5h9EPC2/HjTkcawv6hMqQ
d5D2E8CzG3Puoc4K+wjIajRKFsfz+fHLasBpn6SzP8iQXMSuhpWiK/1pXfab08+Y
cjEx3xNKQJdo2P2g3ywnK3EC2SL9OZxh+ZOv2TE5LL9+J6vWR6+LrrNLbIHC33nw
B8LD1g8g95mc6CCI3UYlEGGPG+pxlJXymWG5tM+uI54m4j8kI+fKAMOBAh7yVjHs
6kNcu1mbf8EEuVO7Rz+tRGMC6NyEEHcYQA50eVebRnUt35yu4y8qFzFATa1n/f8A
XVggK15fxd1CBLD0mr9sh3DYYR5yqczgydvXluJyDl3+r7eh1QRetkFqBlFKEFuQ
J+p7yOr/oRNBQZCcoOjwEY+bGXj6lbPPVW36YP9XWkIXxmhACmyS1Fd9DjTnyGs7
w1KeQXMDTme9zdHQHOxOAFHKL3ZpqGkDNN4LrZwFIFYMGR+/Gkw1L6pvyGeGyxGl
cBltLN4bmwEXj9/9tpxnQYBPfY2xA22LRzFtnMVyCKBeK6ZbdembNbSzfx+xfdKQ
BO8ujfYtQPjeI70Zmx/06eQjSlv74ENd17cbl/cpvsjprVqgQaY6mzVrnLa3P/KG
uPoJbQsG+VfuN5uWuO1A4gKV866qvtYvQTDI/qV6FRejx8ElLEomPTm0zsN+k32+
mhRJN4RqatGBsY6CVt4YebmiuotR1fuJmPWSxCIV/BHi8uiq94iqLkS3A2IJLH64
Yj2kb9Bl8226iQEfKtkeRSxWly51bEimZvd7kUVoe0KucrqXzafMHgaSlDKdiWL9
4hW694hToEcRW5ZuXC8vWs3uFpf++a0G7NKkmjxuA+CScHVBMevp85l2cslBO4xz
pLk8na3zT6oPlZOGuW7ju1lKiPKFA4buHddZRMTO+mrkqKX+9bBAvJA74Wk+sE6u
14dCwct1kn7GUj8RgMChvSurMEC2RcHv6vU5+2VfF/dHv5eNiZSglvclylYGOBey
JAOYkXsHt9emsCAiGnwS8LYXnLP0PxlmYKymXT/GnA8kIT/wY8227CfA5FS2VzLm
kypOyGGeLDEX+6Bv9Wf/OndQBNz5fQA3Ihqufhj08Sz40+N1t22qbd3CguOdKQWJ
6n5JXS9t1Q7/CkqYdlambmMSbUzBMnOapdLYL5UFF/ePghtOohWjYq+Z0QGM2u5u
godJ1VsS09CCWg82o1HhrCiokIQxXVL5h6Stllz6nXdt8H4r72BlvkzwsZMO2fO8
dfbbZe5o09mVs1bAcEYsYTPnKU/HRoSJfl1qtUxVJeIlrbRUH9DH1RpUgAkdONLd
d9YpEIsAWY3nW1k5ycNCFNGEWEX7ziqljrJJisORuOZ/OzDu3nL1UCRLbX+oBRwm
OYMMxCm/yQj5lnqx9eS4hvsgBGxtMM887NLcF+J58h8IwB4lE12fRhb/475YpWwG
NloSUycJlx+lGriy9bgbUDGyPdEh1Xk3+ElKXwkHfPvsO+IozDkKQw0LUM/Fq1vx
MWlS+cjhrA9tkZhiVDl5594EOIT2yAYi6iHpsGKHuF/4MhOtG+JODSrxRoQSjvwk
VhrIEOo7Ba/gjombsB59GYd0ZuJatrfY6vc/t5JjyvdCLf+1zO+qoRMl1pNY9i33
P4AbHrJyGdLcEFaViU7M5RsbSjWk0HHfyVA9Ew1TMlxHogANWi5eMNmXyEXuwKEt
fZQ0NhPCXD09lPADEAeqzDrs1yJRD00iY6IXSI5mHPyndDHwMkk3iwxLMwPgp1R9
gPlwmfjW6pU7hpgOSSPyN7aB1OxXd6Lh7ZQhz49eaRZyIuYDKdDX9qLne9M82d+I
MIfBeqZZRrUtei5o7q/KpvqVFpSA54juWBcsfkWHwGKIYV3p9Vv/iBQkbIY1y8HU
d9mRVu26JHfRKP5vC8+IDOYJ2wAfiIzhDsPw0/eDGPO8aTp0tr4myTuiRu6+qq+4
hXbITvSefHiro86jsK6SRRPY+RlS+LefYyzwgz4qNKKZ6YmGm+FH2KFQYkNA2PyP
H0NyaIbtye68pMem5e5w+8w+ZZkXFejJr5T51o4BNSTEgsag67VxjH+Y9T1Mab7+
LwrerNxzqdoyi1zZxzLdPocsUzFALLBW4Fa8n3osf93dhPd2BOZBIveihbzRdEgE
JxZyFAp7jk96eMc+3a+adBfCfOQQy7uyVBRbx49IKfyGxJ6gMmsPHLVJQKLlPiFg
PaSOeAq7Ufb51iUYVQO/dkGex/iMueyHi8gfxkwro7qfubSYKwNrNo6RaTOtgfOm
DmCHg6YYulTPq8s716RFTIGxTkPWXldQBGEQMdm7KcfUCJXiqz02funF67MggCxM
4KqL08H6J3J01xZFqvqbFuUyWoN2TooEP/52KOaZitBt8FtrHsslEQNfHhpJaGV7
kfo5ISd/AoL7g24U8icymIvtv+dsXFhgesfHVSJVGfUWt4RvcBI4HmMGbm9LOGLs
5msj+zrhPSoB83E0pfwcsjqVGsc+xJttifZ0g8Q9evD/XY0d0ap2FLkkJ4EAsVXs
AaneqnCWXC0c9ey8HFvR1Nv2h1XO9+tejmut1c0Dl5Jgo2AaPsRpXm9dHONCLj6s
l4Td9zPWq9XgWYeW4arLcAjpmAUDs1LZPMe9opRSs9pUslTFNVOnhfGyQ5++/iZH
PBHq6h/lfC7YHKd6S+G2cA64uCwJFCsVsbvrVW/xSUsuW5x5Kzjw9Id2up98acl7
5EXEAdPbp1djWvEgoNo2ghxwMkK+SoJBJlXiawmJHonKfGoAd0jX6dlC+TgSctF+
ho/FRc2cvKdB9u0X9Ot//XUnxglJuQ1+IPrfjLEcUxfrDUyd9cIHdl72pnJMhtP6
lW5MnDD127XANLLZ9TvfjEhZXoSqwmcyxjPEKkboglCKZb6PeXkA8q1ceO5G6cGZ
Xt6//gXztHivaLzFMbgqPiAPNIroIk9nuBcAwlakSLCyglFCk50ytWIemUTv1dbl
oyOK2kHyo7ChDfvlYyCq2XFcNLahAuy5WYIk8m3kcannU1V3J5XgdESoEMjZn6lG
56EkEAMVHKYwSmBzBkg8fo21S0YbaL3qSKnNJCiKgPMJW401gK+Jg2Y/eeBFnk16
LPrlXPKHvhAgSwQZYQAtTROY81Oo8M4BdC/qwz2W9QQIUu8S3rRDOy4QOh7e362W
LfZ2Px11EKc2xoRgtgnpa17//efAvi6nwSFrp9dfmx7g1HNt+UFba8oK91iqa9kj
tkycV6ahZFfC2txaN/Txe7mV+EK0x8v9AzfIr8dcFYRv86kKz9mcW/nivUd3KRCc
PbsRUwDx7rWuxRmNWeEtE6e1NFiMul4CB2bISlwbIegxMeBzn5zySWfwQlnvUG5k
ovjPisC0DBL2O6C0/zKLee8UUfPPA+kZ3VQLJDVk07o8uplAmm9bBrK/djDBQTLI
dUkVfN1U33NUUsOh3tQqgjWT4T19gjsFjJIRZevktmLbQPLMldyZf4JK00APlnlu
MEcjLM9vb8kNINhfSNVBs9101MZLVtr2O7CVpJ+wgWqBtz/PoGsXBcdBRHahz3FO
ynbjs7yrAwgaiytrA2+Wa5CmNa1Stk25XM9om0iRbfeO+lulp9q4vXDRRTRkwuH2
UJkCWClDDqE+2ZH2peIr6EuQ1BqBAap/2uQwCQwWAKpPvOG2x0Fgm60rsKY/X6k0
CGGXLL3aQ3oWlMNB555YpcXiJRYraRwYb1yP84hGhmKRxNRV64aL2Hvt/IdHBkIl
fGR9FjnO5QpNqtyjFieFXOXP+8nnjTN1gUGZf3ruzwSdZSRmE4GUsKIQdks/Klnu
gsRt/djNLe6N1ck36WHwTt3pJDhGIPgRZogWWoKFb+6q1e4w7CnrF0MhGt4CyZRz
kQMhUl9iwE78LXqNNkU6XMynY2f3uUi081FnqMtWPt3fCshtxZb+QnnteEX1we1I
7kgJIaKfTOnTDJ1YnRroQWzdU9ZtfABRaDMFQeI8nXheiArzzc10D5QtPbV3fyAd
bQz/7mPAn3+uKUVHdp8P3+Ouw9BNUuoi0KVEfHExkPok0+ry96tvREzj+1+SOH+N
LSGRjwd73G/vDtexD7vv9jJOy3fJ8VVBJhCyrXNniUFxZbf+PpGatuvZQPlFgXgG
Y1nIZJf2GmQLN9snfNdq4l/KGMTYR4QaA6zyM3fQsWXgxbPo/k7d7jhPTjE0k84i
30qsTPtV5biPCQFRBNwhkWVNrlq3GPuCQNctiGhzS2bikrTp2+atLIj92p5uWMG3
/ZEeaCJDC5hulPyuRuCqQAxidmXPNZBrNTRrLVKy7yAvUw+k3GR3sUDJPmQHJVti
mif2o1fnpmwsUafc5Z0zdl0sxdFUr0n/Q+t3/7ebEmIcHXmoXu2EWHAZ4kny7gDW
NfZ2HvXW4zyatyiWXMYjRoDBTlC3OJIp0gir/7C7jm+XqON422Q/wD3qP6ADaXRA
yK7/839IBXva1da+6g1tUD7oy/oPqhc5gnS/mRPm55zHeequYjIt5+gR19z0m4q4
apNiJyJzIcNrONKR/KeIGN8BAX4yQNyVtGe2pwIDkFtU8p17xEGDvrtJV+YMFPv5
G+C2pKHGON7TFI/uldpF0bdK+X032+Dur0a+KGne+NVx+/SgvXUGJfgUob5Rf/iT
exo669LGC201Y9EexyoqoLh/XVjUTeBu37E7donw4aWXkdCxyAbwVVcReLfka3rQ
pi+yN2c0MxyANUqv3xitRZ8E9XZ3ChKChIpXXnwy3vM3sm7wNfNVGu7VDNfT02RS
DD7g1X6X65bXlrrUJ0eeUI6rhlvg3xQP/WODWKOlcL6U3qeUPrGCe2s/JNehzUkG
dkOJ5vxPUevAEo3DPAKIXfEtzPAm28FarfgRoSkBjD8uUXXDvyInfWypWqN6H0ZG
CR2e4cWLvA4JC8xHS2fSUC5suM7npBMU8UrZXRLlhkx34MOxp2Gn4LBoOxOeRR6q
QNqPvabpjoDNrURLKUTIOfJlMDT6OJT1FXYa/zmcdZMn5l+wGWoB5kxRO8e9/f3e
ut6+axe7Fsay/tgTyjS21Qlfbs8fkJFl0EH9/cUVQS+QwBneYqzEUCRYjwXesnqg
+1miCk/8lo8V224UTWRWlhK1sDSa4/uYFIHaMLfBjHHgewys1KQuJD/VFenGJLZ5
m/330FxJDRaJ+e+SwyiWsE1JkwR7zdeLhPNwCdg05sVNsrrFk1H+De2B+LvGji3h
M1VAymp3cvS/Fa7PO8utnjy+oO1KiSMU4BiuOdsaIkQ516NBMa29Iuk6PpMb5kHE
OB/anTjPdPEAeJ7/cAAsKK8aqYCt1VWo47nghOoZKY+1WY9qaGFCphsQpMx7v29d
SOh7K43h8tmZRjDk7pa9uiryv3ONUSpeASnlEKhE1OwLRPzT0HE344gqcRGGScd6
+SnIrMC0RCWEjaYAgsQl0/mjAn3wrA5duwBRoa8ssw8yxu3O+UL+ttqN+/OD5/Z9
tEloVRHXqfZdV/XOr5aIk1iyTuhCkQGYA4ko+uoHkK13E6jvXnd7BWagvSipkFMz
ubmwR2LfqFHWxh+vKJ8fzdC7fBNeII+8q8vwgpwTIWdThc20UW5si1CSZaCENk+J
vsg+sBN2fZCaoX2fZ8Eeoc9MRnoUvDCcbP2QQo0huV1yuEkwJXEl4nlOM/iUBmOM
Tf+Rzs3kqpmgy+T8BgVxItl+OAOY+cpmoqtRnKZicz6ReIjyT4FtFf2vYZdNAHCt
Sq3z2XmaEJCTlhEy2U21qhKFsK8SSZH9px7VWqSomT1PzA04qKwJHH+lHAn45yx4
KEkpLs/X1I9chl062w+1c4aXV5WI5gOJw5YR2M1/TH0JgFnQ9SCDx8FS7lM02hpk
+0LA+HI1LzTRiPpxi3l6A0jUWn0nVkozsxaKaEaj/9NsPDziPT/IzBL/jRU8hQu1
k/6IVtsx4ddyWp5avezvukQ3k+XmLtTJmq7v7+hHuKPe2wMPil6Xpn0R7xlbbWCg
y6sepKPJpUNVI3F7mS8CPeV7aQEPqGZZ1aMHHL7hfxyenOhLGzI1ahEVswnPckhl
Q23L/dCdyE2SgsmIzXnQF8n1zPDpZETNiMflYXsGaKADPfFVK8F87mP+eYkJgZWI
6NJD18IvJG+XWr+hLoAE/jBj5jEsInlpC8YFXs6IDqjaxsGa6acddf/ChvNDIoAl
PvZQAQWSxTPUr8qNQCtxeOes4UwgirJLOcDVH3q4PK5b+KbyONkm9tIpLxIl0LLK
PJb2cU2KvLyVdY1syHOFm5xSUqYpHwcmodSGwVFZgJnB6YXBKLY8v8axNQPmrna3
5XO0T+NX7RzaPRGrLFf45R7KQKBMmFLOuIYRFIl798ovApjE+MDbNWhAnOnbkyHr
W5Tg3wzw7Ql4xMXg9jsiArVSwSQrG3gmgSu73eF7pi4Wph8Gc58v+A75wSy4T3Yq
s/VLHEKzJmrRTVeM+kFEpWUtJtFAaCQml0ckmP6Jc/zVvl0RWlZRX+Or2z/7lbAl
6tgN8zPIrrlTo355wmjkMrR53ld/nPzor9Sf5obUqWQN3VK3GqP/doZ1BRBGjfDW
HLSPAmRW9WmLJTyKJQtw4U36wdF03PKLx3q8bmkZyDbrOE5BR4kl5Vf2JwN/UI4J
2PSMQf0Djm3ELFQoB9Xs6DAS46hoOuWXJiwMERDaCtTz0IWLZW84dd0ABCPQaX9Q
5vmPGgUeXzyfcfOEspcT7eyaS2eNhv1HeCY5na3kFEEbMNSiSDJy+t31r+aOOMR5
SSYavdg9yWzhEwGqHGupOCczTfTaq3b21MLGAYeWsTUkIaK7JSXUR6bD/uvYMftZ
XnDNnAZqVLmY497caT4idPJrRjQhjApr04n3rU0lc272muZ05nqwNFIG9gjHiUd7
t9gJoo3M/AX6dv6VlM3tJxHfVb/Wg0X4e84Y6xrerywP4scKcIKZs6OLtgAlWa12
BXrkwtJhnHI+srBJdPQiWzTYQA4CWVxYyzIshRRO/iR3hSWKmwy+8769rM6dom24
xw0HwazDkLnUEti2aHQteNi94FdzzndfrzCqZVwx6RrG5pHCJjxjqAdUou5AlkpG
7yiBcydI/vCIGT7JSPGNN1CVi8Hu0gNpSyCOrLaF7YwJS59PBc3q+cdj/IHQIOO6
jFYHxr9PlY+2XrJhZSBDaZnUelx5vIEoMUN1khW5LScYGMGHb2WU+sX02Q0mI9ge
CK0+L1/kM6MW5lexU2PwLS3Vp+dbbGiRfSeyzvN4BB87EpIV1NQwsr5oNSzhfGnf
SRYsLL+5S+CqjF+AoP3ZU7HdlGdvxFgKH4P5+zJnmf83o+QV5eGVRgszdx/t+Pv8
WkZWas/rduMjqiDooQ0vuR164MjorcW2WODRIcIqKpGZ3M1NHIBqu66QeQOaLpHA
A3Tz/wJpEYQ1MkHWTO+PuFaAe8fAiS0388YROh69HQ8ZDw7MWaSJy2y9xaPNuD2W
h59YWRDzDLZwEMcmUNnGslaZqHBCp/gYRfDWvf9IgW9f8dqWE46fqEXWZzsJDf6t
vhQ3qJvSP2CAm2uBfUp4vwFh8n/AYBBq/Eh9cut6BiebBbidEnjbqBpIs6BqUjSd
l3pXIrznxXfLhG+TeRqU0s53D4dr6NP7Pt8YsCyj3CdktEQYPkLtZvZrKg/bi/Wm
OWfp+nrDMnOKjE3c1ld52N+RXZWX90krGQA2Zf6az3kTKNGnfyMDq6BeS/TDwDrF
xqpshUfydBwwslulzyHhsPanl1rV58H+3Mz0+U1klxFKqeXTN/ZPIIFjYtTBExHv
HEa51f5BV8JbRLrLF7yqTFhSqNVw/zJgYn3nfqze99apmrWo3EmhWwFq9fkKw8un
dhLGApU2iAn8xmQEV8WBdYHLYaPwhz6X1iUVs2brQg67Km6POJaaCl5DIgRbLC+C
WHFO4+t0RCks0vJWwmfrhAUUlrXIusPIbCw7qA2oYxG4+dJm1n6tIrBd9PvxYwla
W5Q/tty+6PBQPtXIt/w/acNGd791LmPVn9ezRA0X5ngEBUi3gR8DYf3MeTKY6mYd
BlYQMpGeibq7kNrHiOo8Q8OcOfsavnv7nq0jslC3convj1s5dFMJ5nk10Xz+DJpo
mO2qgsNeC2pMsUKEDAqUHjlJ2I2r7+DVEPPS5JdWZFexcs5bbMjoRQD8bI3s54Wa
jTxV9VhxhrUzB3On4b0alKsyX3QSHgBMyOnP8o7n0eXLl9pkUPT1CYMaHmuwCsNS
x5//WmNwEiQkVdVaY23H+EyYBxhs/A6EilYiP4/nK3BV/T9ytsdUwJMOP8JBvguX
JHbVHUTK4iyD8oiFeVfKcNiTUHq5vq3N3V8LR24UDMY/tf8Nv9PbKvaGiYG21eo5
JNw+kkHnB0pWM/R9Z/dnw30Any+l8NTJgntB6tGBu+AePc4o8vgqmpODtkWxTkPY
IXWmwtaGiD3gTUmCnA3caD4IeyiX+PCHeh/2AqfFsIusWSWPUTMkXGUbXBsNX5AV
n/9zsBwHNaLIy+lrAIUOE/aAxdJb0RQ+7xedMioA90cU/BzP1mrZvDjcdACl4X5K
SlE8pVpcgmUOX/uMe1tE4GCbyJnVqexm0ImJvtixbiLVoR+payUeE9koQUGK6XG/
7iTamT1alZnxYcghwZ0SNlki2QSHJs82gBJGB3hTyWJwLr60NCUek1aY5dGeYMsp
4ReGMLwCpyTGN/5b7Sayftdy5GZDCRJKQywltcLFFWoumMQZmMKzNu7OPOXlmfpm
QPpensd1zbKJSQRLnSln54MfBFeF0csWReJdItEp8ykhWJdsPr8N6Bp4xBYBMCI9
gzbQ7sKQiciPvivNSidNAHcDIPFeiPas0s31EA1Zh66CUgG//x+KmysIzishOKDR
2JY+Uw6u8Zis4/viWabCO2yFkehpKJq28wV+rWrXZnDGm0VXLaAXXXK/s2nNHzmM
H1IvpK/r7AW66uDxiiDM9FzrLl5EbHc39vSvoKAIX5nRJOEU5BIN2qEyinbl+y98
5HRiskRI0hVgK61/PhgU2IldYJTe6/Bny9bp33peDCEIUAh9RdHdmd4mnZoK0rqp
yuVtUaZkAoJm6PyMZURNugK1uL1Tmv4EG8H22hTuFpEILVBJ50msfB2sG/xIWY1Y
B8z0YjczmtiF6rX3xLap5WYIaPYKEkw9SZpEHRbnrm+fjqk4tecZYgHoNNbu0OEA
7EIqK5n239OlEzghgIyzFaZ89h6f+6fyn7F4h4eB7O7ZmXGPzqFrXHVAq0la2zKz
TwvcynhH77lAxAVMv44hUqJm+BjV1kquyGGFcz6G6IESkY0dpWyKClE9NYt5/zAv
aZEM9HIF+P26pJbNaEsOPBOcyOzTURQ8Fxq+DBxfGERzFZ1CspuaNNVDpBF/78Pk
yvtMVXbtNzDFOyXxafNvHKwdZ6oXasJAEVHcWDBnoCARG0aovfBVkFVBlnkTRhFe
lQdNNIAj7T3qqU5pkVYRjdB9DOqUJ2IKWh8Z9OYMud1oXnMZJJIDdbjfUkc/fof4
QkwPpdvWAf0dcLM9f2avnBmSBQPTB9KkEcr+nrp+QfwLnoH/NAc64DMNNkHdCoo9
rOnE8sk0MxgoGXAUCOSPAF7/xEoXCDI5GemHFfa686M4NGoy+GFs26Ltu+tHWcpy
749rE6hN5y6VQl0Md4e0h5yVvsQtMoJGn/oRuzko80+k02Q84j7QuuZwELnrORbl
vTiex8FDDlpTLud0pqxny8GD9e2GRVPiTZPOaUboeXnuwLCMBqqDloB4txNPJ5+t
Zpz4s5xS2jJrC6L2QqgP8DkXsj61/2gNsVoY6WhIa+FecLIxyDw5ITbm/s66GRDg
uLprBpYKXu+Dr7YV+Sxyp1GcCeFARgqB3S3CzUCRHujaQh7UiH4GOoAPSdL0YEBS
ZAGzSdx4IMgnIAg6z9eduqkXpy2N8NtoDByCIsKiJWnM6RN7dH1EQTjAWVKftn6n
/saSYmjUNHxDNuaVBP8fTtMh3NMhX8xfCLANNCfGONlPDCwr/4M0wHAia5WJ9EzX
r+vHEajwrHDh270oGVvBQfawloGJnWMyrFfsH0B9BJsoUzNUI9vI/UGGO30NbHNM
jBb9R21k06FefGg7QjE/gprzvFr+bZbA+Qc1Pa7dimXB0lhd/XtGd5Xr2es44hNy
MdPdw5/MZ5n3dzbHWedk71QKc5Rkhap8TaGeVXlpM17BzJIs7NQ2kSynGLqsPA5M
Cyr/Nm4R/ixZrwNNPGBmGyA+GxpiB2alP47gjQ695YTof+glp8aCuWu3IDzWRHr7
q1OObcvAXmgmw4jWB0sMwXF0PLR3Gqlxd8X90XX5uDUrVLbnLfg2ghh6g6qU+5xQ
MsCD7PAOOXPcIxN09vdfHF0suCKWUI2coAyDh75B36zhuteiEeSd61ISwqpCTd0m
wULKVekudpQOCDozXa7IcNHJArfpQhqZdI6qL4DzTninoIysrU5Zm5ZB+jdfkEub
/iV9CzdxWreA/aI3OOVYcRhb9iX9bLY5XPZgekIVBoD40ZDhvr+FzBf6XHv88REE
9Sla+sEM27yMgfvFOolK3/74u5vCXBm+Jt0i4uS4/55Ln7sJvUG5EsScqmq2/XRz
nJ19sb/BJDNgY1tEsQDguCTP05bDNf4SOF8TTfbGBok0kQq7nvkJGBxyZesi8HGm
4JfKCHvyUKGPKnHxI9lwsNbLzleSD1W3WTxDkCI06pinXPdA+v+PxVX5b0DIC/mg
2r6T76vOOJl9n943bn8DhvUVPi/06t8WMtCX7rZL+it2zTgKQTqfROMHDE4+tyzj
WDrJ+iP7SoDBxIpmPiI73pnDKkMThv7OGlCPA/80dJPSRoyi5iwuy48raahb8jIK
JdQ4ib+y7wCPvr0nBhdt9b7YojxmzwhOZTH0GUmXhyR8yI7nsWzS2WpUMCad7Djh
5sHPfO29JeHUjWtOGebxM9W/VDbKpW8na9Zpld/LBsurjmCAE5fI/3/apHFjaGvn
o5x/X/KMtQgQHcZA+hFQ2We0DBTY5l3tf6wqzprB2kBKobs0vg5miQf5SXqZBozX
WD6vDShW/bMOBQd0sZR+fvrMO5aSNPW+QBzrZBIR3RbF9a66/izAocLcvHLuirVw
PdvzBFFbG6MEhQ6yXlnKyvH7VhDVHhY5Z3nr8++aK9SRwXeBnfrQfomE2MU7DTzV
FfR83106NCBefhmBvKblaqHz71qeeKpRoJuq3K4sAkPdI5ZiT8/yhdxjxq5Uc6sv
SVdMJUU8T0mJT8WfWPZW7V/YV9IUhkrrJKmL0YJfFRPGPz0PK23SUrYevA1cxEsU
lmfvnMUV08O0v97Df9Oe0x6xlfZfV9NXM/nxPPl1oGnm4M41A4AJDNzKh7rZ9g0Z
ZPZT1DCzSsyZI5kc1HdJ5eCyLYyWK+TWlL2F3rVu33TUjSQF+NQgP81YOXq1zjX0
VN5Xvi8UDFl7aUFbfq+dJqqtAVJWlSHvObNl1bAa+pe2QNj7SXOdIAm6jq9dIF67
ewwSfbUCGeQ6BrbeQKL//ebxP0MZUnumZYssLgEZf+hozREaETbVgoWZXho0+1tH
to/JZvyKDW+nMRgY5QThS0Sp1IUT9eLI6Gi3U3pppQI+4mIA3eGX0W6EEOfBAfiQ
R8H8TW/T7soI2u7Xji9r5PsU56JRHt0y5CFD8LxENVrKchi4kJXF1eEYhSgFJf/+
QHQojSGeXbT4XXX3fnpQUyb63uuOmiS1QoB9W9FtGuJehrrceS+9zRcFqD92Up7z
seaFQZb30n8LYwRZK5vNgU3QeaRRuhDI/prQGyFqeFuG9g+QF0dT9ug4q8ZT1Tu7
VQfYosO2hHLTZ6AsxPoxJ4+b4jrc3jIucYEs5TWjukbSnr4KStA2X7A1lODTh0jM
KuKZmIRp27rqADcShsBhkeIg263+EBN+SIw/zOTBiWq/FdEHP7TufFhj/C9XNWkG
cw2UtogvvJ4lGJXVWHyMXtCgfgUlC4Gn385M/hVjIv/wX0s/y5ib2vF9Z4bJMbum
IwuZPwrDwn8Bp5lzHpiWY1gKjPy069J5l5t+TEghHweW0vRxboscAzlV660HVeHw
wRr84NTmwBiU74nI/Agr0D2KsrFAq8iZbDTypK4RV6QmdK4G/nRUvoKYBD30zmcZ
lu7pLfHwuRxKekho/Tsku7w0X9XGNtByj5VtEch+B4DwOANecZd5WBgKCuuflcIO
o/ZrSu04YPrbGC6G5w/6x15ToSQFfPQlN/PQvYMOrtWdiAkRM+YPtgk6CxtoY2vF
CgeWnZhxiD/vhcXlYe8CxmWbsn0nt1lR5uCqx/niUFmCdmqkfFg9r1Ojm0zHEXEs
1gZyxDDHdyfFk2gf+S4SV4lEnux0Zf5zuxawMHYguK8OmKfJG/ZtYVwXF3bv4WCa
Hs5P7Uw+ZJD4IoZ43zxmh69cmq22uHeae+UsR7UPycpnIBqaLTSjbyEvHqGRsRua
VAp4Wv9Lp8b/kPadSGrEJXTkyKgYGuuV2IxBwUACxDDyPOGsbkK0/AQA4S2IHh2b
rlYMsUYyYbQ4BBK0xSlWHTuScbkbrF0K3kwniDs0V2If6URJLH/WX0/zGh8ZcdEp
MqtCO+i2ew/TbL14AdF6Ep5R48f/1IxW6OXlOiVymxMIRDxRtQqc3tPYpe/ZVDx1
PiPzSDgbdWlCj1iQlAuj3xv+jr5gxTSqa0ER0ekWHM8u8uEew63OkuGGYrV3VD9M
ooFuS9P/n7murY9SuqzYdr95Mjflw/dcvXT26bedGNulSvOmfz65qvAWJ2LFYZ5r
IO6EaCA4Gk3+Si25JGg/YA+JYOFpeH/rWVI6kQPtcL1AwnH7dnA7geR6yRmsRQ4y
u27TnsPHF34jQl68fua2D5LU9z2ejotG+V+ePr3J1ao7njTFsC+BtKBHQJnFvdgS
nGVLMEvSA1Rmh8zJd2KW9x2L7nJB3nU3qxWBjg5Q6lDBf1TBxKFzdZdL6CIxTeDF
3G03kKNYERN9gEhp4b1jYhBoSBw8HnNRFvnPJZRH4B3FU10/m08REpahpc5mJ9Ax
DP7BVQFK90JXky/j4HMto3tN5yxHlXlxiQxpq5MTOiC7bGlqwVYGG6WfVQohu9QQ
iI1WBFosWLvprJZd5oZ8n8XNrravRAFI2ziP3zGK3WL6urt1OIi6+eapIEM5nHJO
FXs9A6g8BiRlgHLONaK9uR0AUMpTrpZ4D8Xyg9QGUDoymN0VqayckWyTfK3uHrwL
fBVTtqw2eP6fVXaPwl5uRhUZMRZyCG05JhIGfhIhXs63w3FrHFh28yMFonCk9alI
sbTQr/G+UqtfLLedhr284ngYT50THYXei21F0ax6AgQ0fzr2+lnIQI2RRo6anYDZ
tyuteuBGzkuggVBJqxToNC2cYD+xH5aPtjnY1Mf8hlM3nIf2EEfdf5vTFN5RV6km
u10+NeDDJ0x3C5DZ4CKlhHgoMaDVY48TaD8zVBVPVN6900BVKLcQ9g5YNioKKvOn
AXrPC5e9TzKM4YjYHpLNoAuWpviGfJJxdno4urtBk8G2SZH0V29vsXvT3mjThRmU
HjJ/PwwJRQsCs494SjK5MDw/l3bukkpp9r/ErBqRqBitkUv2OAtqPqk9QOhxrphe
BYxF6BKHKyM1wysyPinP1uAL426EatrfVnmY/m3WaS+pZN6MjJCCU5vXR7s4nO42
2z2cHsuidg3pD8KUTaa4VYspcSW6+WnPQla2yKL8FQDgbfFIsHGqubpMX8pc3B8L
mZBl63uVXTnKeJrcNt8B1xzGalBEhi7hNNvV1uDp0YCBjZVBpR/8EFMMfcIIDLjq
/YubXWjgGnU7Hsg9bjfZozCT2SDcdTCmap6rJIVxxgCwYSEQgIu/HYTvKnaM8Ajm
aMluEFP5sRH1MGZwqwCWqgxgBDILF1+zR9HE2xxCrcSrNLaOAi/Dz50GtjoQ0tYw
DHwfQtouW7LKwdr+0QtgYvrivXPAzDIexPhN5EJaNFUpsa/vVhEjKVy0BFls+Rl4
BOwn6Qf7UR+a3dY3wh5TlR2761eOJX9Adxsi8NGaJS/5HEdXLYtl+SEdm6xglwdL
gFHskR8bd5RkRvYSMD6asvr3aEYF/sTHLXIJSHS8/XlwlJUbw3vPsryIKOQ5DQ4e
ZYnM5yVLNscrZOmaJH1ZLk8yDHCxG3KM4Hdkbys46tRgUQJ4YBmsvSxv5Eb3zVee
DxzLQF11ob9tSFIhYHPDT+dDAlydHV2csS4RzvJaKrTtyL+c76S5sxb/eQK6yt4V
y5Mt5S9DpuViUupcIgXAGPAeCPgOe0TO+qNAy30v1KV/CqLlGV/fmMOuVQobJCKo
BLJuj5MJOiHo5oZi6wsIkFQcB+mFihItb/unghbR0cENnIvv0T7u8towP5VU/jqj
eX9zomYsPySgnPvMO7vZWCpZ9cAmrjcAjqtzMbKwWNciU5NdKJJJAQF4f0AQyECh
TcjBvq7QRyFL3Fei943iCGoBR5HJ6uvCuXsZ89q3t+4gDhfgTlhH47IKRE9x0Rt2
B/RzeGxCLr/aWwXe4P4Hy1gKiYg+DAL/u/YCYikIJjNGWhdFkK0qJN53D9Vw0sgV
IQrdxKW87c3SKnjti20FpX7QG39BwkU3yjbCycxk6FsSCi4ltTyQnfwHgldUujPs
I6ZkjjGqvxIXWBB8CkvWSkse03x1cjv6qqBZey3JJeqsBO6Q0rvSRpLv4/aJuxHy
8nUqKktRH6UAwWTLZQzQbmV2Ry6uVraBgOxeSO/wZ/8xjq4F32JHzE8mBne/XYrJ
VC+tzgl3NDag1f+n7RPL9MVCLxQ3ti02Jcoc7gGhHAtTx8eTL8/v8UNeKalIHm0f
MBIu2h3SCbo2daWQB1Kw5d2Lm7Z1mmKqOcOUVxCEQpQK/5Yq/dNO/mnPXq95J+Xz
ZAdN20hmDcsbC48C2jI4aRlXdll1sipziVq+JYE14GtPUpzWhyRI8+lHVljc8B50
ChvfkLajM/dkaPUdbnFUsH1NRsQ9VEyG7eM9eOM/KV3Ugk6SO9A90vnpBder3GhH
bORbOgkLbWZOl9J+GIYaSbjqMP4j0fLh1h8i5R4+EdQlcXGBr253eiwc/0S/qXrD
803fYDiiOqkclSgXDsMG4HYd9E9YrOPTk0jjHQy5Mc8aeARJmcQoqtx+Z1LXJh5/
IzuZWMEkefRZ+OK8x4X2jB+AMpc5cN2xllodzVW0ocmElaDfO9mjgtLCUStw9fXq
vVZvh/LOxCJ7msmA+kJpLjlucmcjCr/lhl/x2LK6nlQ4+bBqZvRA/lZlCTkmnsdU
MS/n8rSiRTqJ/c74fFzCwm4aAXZeWFOWm7mo6wWEpbILwM3YyuxdIErxzTrmxh+2
FTLxMTubEE0Vm9J0VAsZ1N7aB7401qht7PzM7/CNcbnnXIrZRCzneO2NzROhxFgP
IvYBhZoS1kQfPcecL4aKMiYtKQA+kG1dpYHUX7tN4+z8hNdFop+c0eXH5e4ng9Ga
EgWqEuvgY6EUR2G6+fW2+AU6giFXiyEA5JDpHYOso9vIQR0sPNDoeyl744owx9Wz
yrHLBdOrj1w4XUEbXY2UWSn7IgXCYigrFsXbpWpaoS+lXy9OVhmVdrivPPi2Fit8
lD21n+bDJua9mkd8pZZfgMr51CISUJdhjyUJW+NbEiyxQqK74/DYTVhtRXoi/CEs
7GSNO+vBsqGPD7Jf9aN+ILwuy6dxttm5VCiSIjcpiMrrg///fNuWe2HWdcDvUE29
PiKX/rRoC/JiZijuZBryWryNiPhrNzVvegBn8we5xz9hUGhqQIFKWw/2LpU8zZwy
kaveXQCD1lVvLnOvkGWMBQDX+uEDtBmb+8bZhqMRVIvmDShrTG8P2FgIysco0yWh
io2g5V2Wt0zOlc8dAt/dz2sjwFPbsjNUVDXLDVJOhFxkveC4DleUjCB/9tcwonNA
NmGVbBFRDBRaqF5IqIRAFqZI9F54+A4AaNC86ctF+TRZPjrNYEuyCrU/Xq0rBqVm
k1EUcILiiU/IluVxBVe9W+SXUGrYWYMK8k/oRZ46ZlJNgIL7iWB3EaW3oM9SUQnW
Fqejq1StQoZe75Sl/hgRCGsApqGUFLa/hEhE4651sqWcjdzUaqPz7OzZxUxnDmhb
5WXRe/+A6C94f++kDxNunDLjO7CLsbx9cPoRHsBVXx5qeZP0OPD+HXQq64ffzqLO
9Cdn7JxHTdnn8GCsjUoJ0SEnrZnbGTgqcfBwz02sWrRYcbEWLmyWxOHuFSa7rK/Q
r6pqR3RiSyjv52+psBAZClo3iJM/IYhEv+Aawq4MXD/TKCA6lGo6WCQlObW7yNtt
BUDqmE946zwDvYF06/Zzjqv3yYj2Rw4s9ryE0zK1q3REu85UWVysyqFJu6Ef0CgM
W0l01gfLUknMAf2Uv+ktSu/XaleJWLAn91Z8UCclXGL05gu3gcV9ilTC/AmDIWxn
zoQe0SRGazKMO9l2QqmJN/vS8JcyGSPYUhk9GiaxVX8B20qoz5/eGQKInlhmJs0e
wmOsdFw2LEZjqkA+UH74o6XLuTZNA8izwekjn/iihcIEh1flmeM6+lFuDOr+K7Iy
OKl+ltr9UGxsRKFMOTd9URWoWPl4aJLJ1sg+5H4XdkmZUdk12NSgYt0V8ezER1BA
atQzqiULrsGwmDzXaf19Tb5xffn5r3yhyLH9k6Pbop5Ce9xLraUvht2gSloOi0Sm
/KGUE6lUM3cnOu6hPYQYdfzK7mw5cE5beZbkGCbCECGjSz+4cih+OB7GHf7OhRNe
BqT4HqOsz6FBAT74LpzRVnsgFJKILRMRmLraVb8s4q71yg0WRNhMY/w8pgCQWSl5
IffMoCbZK6/mhVzZaTAFwyDO90Fdp+7w2+7u0/fHipD0UvzeWwQzzx149GFKHgbt
5SQUlQnEIvlberXqFmfu2yqutqBoNoyYiZ/Tb/iZAhBjNrlatXD9cePpW4M8zk5t
vPebAG6v3Aw5nwBuL7HVdTF+4qkoPo7ecOeuvBAAaRJ2ioX5RluaX2EOM5L1y+Vj
lJOOQzbodg+m8XOAhhhv0lw48B98caHG2G2pG+PBwYUNKOnszUk0eFdLFA4qJP4L
dDyXxhSv6oo4MaN54AbClRalM0sqvL8ERd0O+ZAWZSjMqW/a0qDnIdNiGqx3Bi2I
vzDoeAiyw9GHEjSJfKCi+LlvnXpkU/6ebgthFcQdhu+PJuWHeyYi9eExQOqJlz+o
75fz7+Vyf4ErEjIgFibjbOkB9C2cbY3fQiNRzz++Or7BlPSZVWSnTUv2/pnguvJf
tvMEROqae2Z1mFHlNQZcemeF2UgGt/U4TfwzW1pwTX47WnYOyk1uNBfhwEGo1SGk
LwEgtVLmFneTDhsJRJjpLaPo/Mb8hWmFdiMuArdCK3v1PpspNmpUu32ZtBvYWlOA
1sJfc8M42wbBvWeGzjlf4iD5ya3SMuWIXORQ1zMBmcPwMxhIxUWVsNzrXuWEApP6
eVmxYqd9RDFDbcqzrTQgnjivp89z5H28z+LTgcWJ1pnfRZni5/WN20jBsoRaYAHz
S3B+fbwhGTvVBIpnYjR3QvZcvfilS3BfIKv7v0qHRgLzSiIHWuq8u32v/HtalmWx
WB/h4PdqPioCrj+RhzEi0waZl2gF+0J2Cnov/oQWtuaUyQOHbtRlQFBWOMkPe4Sa
dhn8vq71Kf3my9hGx93bJH+39UBiOgIIiHSZvERsyMEC4/10aVaeaSMqG06NOv5a
uU2H6XqNL7WEK0NIfz3ApvSGMfwJw24gXgqBHjAeMMy+WQR9+3UkjUU6loO4HHUe
lngn75hNrMzeQ0/fA/CErOXn9JWty+jNY3rHxvCDsdTO6hsqspYAkp05iGoTPUfy
IGHVJ9loFxCgmFhgTqw0d7d6UQP5lxMwkHEWLOVXQxBAmr/+pVTRcNT7V8BYc8OA
bzjuAnpGMSyuytzUh9leYppskMhJ+H0hWMj8CEvrHcnPKJPkL6wjK7wUeCSF83t+
2HW+w7nG9hGBtmWImR7Ipms6ji7EU4RU1nVK3KUE54z884XM5uy6Ade1luxXx0Bu
dJC0uf6fstZEIfi9H3yTe0z6mxv80IJrnq9cXtFL1P0ECgYVqbe2ow6O9i9Ax38j
gbBATWEKnq1V7+4BTK75cepddTYAW83yw750o6Wsn1JNCRhM4UN/UiYa7ahUfxYS
ZIujoDngnmBmPf1fHg21SyepqNG4SAkni+WSYnJkUW92iqXJPLB/2TGAQzQYmB3b
C0Y1Ju5PEgUJr7f/qbfkQPeoGyKd9G38Jy/d8gVVXpsNLic46pmR319BS8Sg5f3b
uD8xXUknMlC3eKED93ggOcUWM0vWOuV+latpmQ1ItQ41p2hwIIpY+9U1tAZ/8Y5m
uhyBAQHUGuaDeSVYgKzzWG2dJ7fR4ZH28Bq/EfhM+vPH6aT7HN5pj/208RHbcIhe
1TyJpzqJtAniRpV01JklrhDaCnlUaZeWzgTLW2Bg2GIWBLiwIWMJC/dGcAXNDBXD
CqUF3HfrGHNa2zg0rqLCHtivr4mPZK4uUNb3yETvYoXWj/Tz5FrgGYHlkoM/aW9o
8sg04rscetkLYfTAIOVUlqW3cZCmfljIQAY4HL/7aktUhVioKWsRP1zSWUemqukK
xeLNG2/taQ8HW7yHKA4+2tw4FI+xi8K/WaSgdFFH5aq2gkiFCcMkInvi6HUUDx5s
gkJU0DOFjN/MCChvI+vDc6INiev4rUMhgC5Wa8gtfl8dNN60SNyuoSmDU13/yoWW
geE1wzMIm/cLrEu62mX75se9O50ZAhDrMmohgXQrtKzUwN80Gtq4nJghxr1YAOPy
UBS2RUmjWEJHenAU4Z1osg+TOu9jyLeRP1vT5hss0rB+KfO69x18qqWh3iE8Mr98
bAWxtXko4/NCKv2zYHx2ziP06pAm3+07/YUzU53/6Fvxbu3wndnU50kWxmix2t9I
2CXRC9BAdvRMdZSMAtKV3uBDtiSzZ7kBl7r445F/1ZMRFdPOpQ40MFdSoE7f00AQ
el8nVD5IaUhlX9C+CEKyM+jU42QLaG9fyRKX4iqNALFP4/vFu5H6ZHJVNLB+xT86
4qdRvellgKezpBRqTbL4lJ8TypPm/dKulKbV+SegTUqxySHryR0BL9KDWNVZZXBj
pWYMAjX6rUGU1qkuFGM9XoLUYJv+nrx7Q9rmiFZb9YR7HAoDy67gO/OiHqFPHARQ
oVuolB/TV7cDqtTfycIpxoVNyX4tRvoUi9SDw73M1DnoHhC9imTaed9fJ5LuH31b
LHEnBX0WzWRBcITDMEg0/i27WezEpERg30A0iQ4wCbnOILASStY5R/i0uQYzGzBX
mAidsg8c4qB9TLdPLyHVx+Vre9t4kb2zG/GVXyrLPd5pnaCEHS9fveJ0wk2ImWoU
2GG6HlGa2oOtqh05OEDTU5eYNjiDAW1vd3IfqRWggnAVOr+DedKrcNrIUI9nONY3
T13mqLwOn6MrRPU/FHgH9mdzXfmzO/1oylC9qH/zFvMf0sr7J9x3ukbVYKg6DcGm
z13rzS2k398e5769ayFotY0U8ofDnsvqj27Ae7hMbjsenqRltAY5zYGgs/kF5hE9
P/9eg7JWby4GDFFR1tBreahuFe1nOk2u2K0P9BJTqwwEzGtpXzs0i1qhSiDIP1M7
SpHv7AGH13XOCrjBamKCN8AUP75ihWtFNnZG5zjIa6RcUSSlBBlPp39f1SERLqTB
O6wRxihBVwdkAyBK7DIc+nLSDqf+fjYtz8TmaRraNvoCPFdUBJK6wrKavhIG9Awo
NDY3xEv5Fs83tWvI2rbtEbrMu2TMKuKZ6xjpd+JOhe6P/tcLwZLMKLKkqiJvtF8C
5qWJ6Ce5kFRLJ5HEWPey76fK+I1OQByg6Hn/k0IWC4kAvAKmEaDgW5KjcsO/og2E
RBuX9OgY6EyTl2HoaLWkFayph8K7PgW05/XcztKym/78j8JPiKwynL008DkegZZ8
aqhR71duWY9gGigTD83pJYAG/xsvXx+tYhgmE4oOY3Mj0+9Z4fs25/CyB2FAeiY2
50bNYgzbECPfFxSMBhKsIkbMHJD7UKzwQitDCNloesNmR5rFU4+LUE19pRcJiZlD
tgYsJZwNSDcXfIRYA7pG6MFmy90UAe2Dbqg9XWThQzdc6GWruN1BLEfHVe5QmSsE
Q4IsK6JD/w+R0fAj7KGGVb75DwKxqyNZ2bC3IKm0tRTXuHj3D3IpxPPthOsd+pVe
woP1GneDqt+YUqHNsu0W/j9EYseXGCeOuolesG97l3b1ZSN3h9kMLdidqnT0Tuok
kErmzJMMQU4s85jq/OU44HtWjZzs7x+XoBkTJRSNGv92oaGLUCv/crK3eNQMV9gQ
EoYAULcjGSBh7aRcE16YobRbjiF8cHay3x3so3FGicjzGszCl8CZy2Q1oa1Eq5SH
s2QiY1rUyecJw1XHUDPQLMrttPU2DVGectBGLgtRNDxQM2Q6NX3kXgrVPCz5Wtjm
zt45l/CboGsATQlL0gFzMItGTbxDSduLXrqr70xg2FUT8AP7SrevzpgRzB5dHi8a
DIsOZzWzFrroWy3NKQmTIQHfaSxh27m9PxkgAQxK9nFmKdZo3ge6RWDHjjIzCp/H
93TJXgJNtbkCkN8tF2gjzWTyLmu1R4rh+juCnZ29PF5uXDGLKpqcoJc02KUV9mz8
Y60m9s5BaAZPMQG+JTolUzzcKeZ+8B2sivYG61lHFXf1urisv6+hT3k84fA3bWmV
RkYqCiGE35+W0gWWTHUNJNKHsdxKbKCEgaSlUo7x61l+44O3Jp3nmso1boPgZ2NA
SkRAJMoeajKW5DV/oEuvkDWQ5FjF8tQN3shDB4NxUnk3uYXr+MTwei0MhYjyknhJ
e0Wgl9YjfCX2O5HUzUSK24hwwJ+B1uXkvOPr199Avk+e3qsTGAcWp1YawGjl9wJ5
9lWugxdUxb1WdTqPSdK6rxYmvZ9m1F5MIMW5a2fYnarCX2LriRF60NFvRKlJoDmo
kyXxKGyMCTNIfHDfB8qbnEHMzUkY6nkXvDCqnOdwiSYrBHakn2T1d1NakofLCIUv
FuIeFDth/wwJhD6dWMW4HfbP1AS3OTLQHYkDlcWF5dsIZKs93TsUaxIyRg9qLObR
41SlCpt1RMdDWz3feSs9vHu8EEgRe0tF0xMKXRjkFK2K0l/z6isCZlh7MB2i6qiS
yNgDh7yo6fh4HMOEpOvcMyp/AawjEmL7EOLzkjXxZD0CI56WAETV1UwPPdMcokqs
B2cQhIX7KecEOGgumtdr2OwsFvlAmOjZwH7xnKYb48T1sTi34T9UrwUPLovDo71V
gDob3Ky4eCz83EHv4rOH7yYsc6NP0YtF0M95L4x5ljJwBRwtR9GwMlFk8SF6INUR
ZK/ckcCEz3rXp6dHD1SzTJXYYFZNC20QujY2AKmWSRdqui2q+leDK61z2K9U9yXt
yToRyZJ0Jrzz3fxiO9mqzU301YlGs0pb0cH+wSHg/0+6QXt3Z3eLA21aUgzDgLD1
seqfY1mhmxwZOd1bZKVJfliRP70qwxrktZJZ7vDuDHObggebIKUgUEVLLkRymOJc
ULdDzKAikpM9X6ETIM+8FcpxAsX1DDAksN/Th0X0fPCYj3+ZEtx34zvP5geAa2MY
zgjaznXYIbQhj+8UGkImDKs1UKaiyB/ATsQlTEOVuXLSb5xv7tc5Vbp4JqJnmmjo
ZdW6AE8WgVwjGgj205unLo0SB/5nTCBl6HSfHTEn0z8HEcpyyLZQx7aj9gd5eIv6
ikk7FpdVi/mZLwW+ZS/sheKah8Xf3RUY+Tze88mJ+bJ+GSZLN9lSPMCXtR3kSWDk
YEdYvI2zKluL+Cz0AgYHTuhLpIcHkqyEevAXgHvfZmTVP4kw98QvaJrgcslH+ppM
qzK3UBTI6KsmL/AbfZIIYxEUjO8zhHwHnid9kjN8106xMa4+IxLl2E7twFrcufs7
+kdbrC9mMnfLmxCsKUR0moHScVKbq2nIvJrYghcUMYK7XdoUhxF8RKIMhht1/dGZ
wqqT1cTW1OMOSTqjo4mb8DymTopM1n2KNEZaRDV+xjgK5papUoFXtEphr2qw2czu
c3ISxRlN4vLLXwpxvtMqkNgyHh1gKhoMWEIXSMM6yJKsOafzQOKptjZoE/cjDDEc
sXt8BKk+RGVtpf/sjd8YbvKItJGW/8ke8ZncZZWB3n6AKF7kv5uAd1b0fbCdRR7B
u+uF8hMTaj7WhFld2FgGz9wID6n91Y9AwmTKnufOOd1bH61Du8whFEVuzd0RNUKE
68j4S9LJ5mJi6xFFYCZjkyBdPZINaGQHHKMq+zUNfnM0ZjNnrW/LjyYvsMqZ/U9w
vL50w3NggDojv6U+J5ak+t8KvNIS1Z+pPCfuDcMqOEEMt+E6bFfC0QUenlQoIqaE
gssCBln81mdYCFztVuUJN9sM8ffLROkyhpWNwGsSAkTWO6yBbkjsQTxhwZcz9gBS
Db3mfWejI3qGIgM/3dcVhOgxcshQp/z+nkRhCwwTGtFIXlUAjfys/BHpW4jCEQ20
ZXlpV9GgddpfhytUl2CJB+OQi6gdU+qBu/HJ/Z40LBOQSFih0dBrK/fQ2llqgZ5q
BykB2GzDHDzJ6tHjMu4+jyVIdcRdktWuU2lTfzL3Bbf2nNVI4x5o4ZGVIPZf2atz
k9MuEP+6MWspHZ+wOjU9NOYVHpHp0x+pg7hvgIHnXwCYK7KXEkfrAW/D4MU2wIVQ
qza7ldWIhtn2WQ0GCNblnZMdhbFEtnI+eQo3iCaZHDlHrCLKoLrAkYsd9wpdIkt0
6HFsZ7D2opNuCeq2UbIgfGM/7aGNtjtT3Q3r53rJTwsO4d4GAqkMLTTHo7a1+5jn
WP8892GJ4JX6IgXJUz9opy7FGoJ3u+Xv41yRZOJ6fb8uLr3quJoGt4QDyMV5EoL6
bkXrtx3PtdAfI4W70bTk/QWoTq9GN6KXGmopBU/89pnSSg8Bqx5iCInenaFI3dIP
A+IhSUnO4XRlxF4c5U/aVGosJO8/d8o+jwyJt8D8nn3SAm1Vw3d4w9F9w0E18+Al
eLVfVhty/7AOx7eNeinZOKrZaj7lma42fSwOV3+um8ng0HruTewZeQsV/LNWnmUg
iKH9Anl0Z93ygw3VA1vdtS/wdzCstKZio0OsB1e4IHXIMGp8WVxSzRttDEvOlF+U
P3jebT5g6HrBQlClEdZ4ClhncR6ErzGbvTwseUuUVOmCtBbcMRFQc+0TCusEu2ZL
/G7Cbe3GHQSR1LR36Un8/E1i2k0bnqEshBYUOj6BgLBclZ87Zbm40nQIYCQ8hG20
66QXXy5qOSJTuhvmETkOHxSIozaMGTy4o9fLi5MCSwUfeQjlz1OIYyKCW84rjmWm
tzRTF7B/V1IsxJsswNgSAGqKcbCL61pF3L9HQ0U7GkCMi1sCOFGU7D7j88W2jhEQ
0f1bMsGG8Dx4mARoX93AsXK0o4FeoJ9MOJ9RGFWOENlnPxOB9MJTPrlIVbhbOOP9
D2GNpUtBqwHbpdTUlxRhBqEMpHulwTad8PiZab8b9VMehGmSV1st1UVgWRqPuVYo
47aHMZULJ/8uPxu7VUvEvcLLR1B80YqDWF+jRoek2aVYR8bCY/M6GveJTQwV8te2
KBemKJJbyA+PhqVNiXgz9NYUAZOqgjorA+gqFozk0mN7PojqqIXb0uyp0EkVZBMO
Y3sJVG89XPI551ZI4DWJ5IAbwO/awmXwObw0wanuvME25c0mPO1RRTReuzHdc4Q3
gdA60zrzTKJ3R1QjnYdr6TvocFxaagJjS9HM5CztH3e2LjblHK2suksljgwpNdov
RasdUX7hNnwdI2IyFKUg24Vh03xtxR0oPlV3juxBTa8B0tyEj3VGfS7wjcxtXi7b
zBs14tA8rZ3EU1Uh5YqKhsr44Jtpdvl1JnRndDxvdN9qF+gkWFjN0y7/PxIwUQYc
EznKD1DVWGi3KsYOHA2nk8/arxQbD3bSZj+M2fG0kRO8GzFWfDkW5cRk+ENdX2ly
0pWSwmvJIYmMlNApRNt9B0o3VrJskXmVxuZqr0wTeKID8VsUkmQj7KqN9MdpH6Ns
o/SwJ4nHsmmsjgjxN3wwstgF7RZXQt11ugbWIyOuOciB9cy/vHNQBpojnyJ+QwJF
2/FXjOfvXILj4Yj6jMjQOIao25Q1ijx6kkqTOixrBcrXPmh994PvWE3cnOaJ5JBE
cLIqDTpPS4oSCqox7FruW78sKnVDJXd2XI0iN53Jtkwc7iCrfgOh6d2yCubT00/x
gTYmSVr/MZFHWMZyjGw73MvIqDolmlphBphHp5NDD2QIUKG7UspPeAbyP6BQVDpb
R01MsZZd7DU4pHWBGf2i1XVTR/Mraw3wiQnjdnIuWVbvq30MJDAHBnJJN4cinESf
om1y1bfe0AiZQHIo+/ZeuNqQIicDdzMbFdTkWL5N70PNE0RBRoDv8U0E25bgk2hO
Mh9WygzbSzJZv+AkJqjh50Nra5+5zJGrbBYH90SD/RPQ9UM0INXnoKKCv2UOdE9+
oTqbAw3O4r+SUvYl8OYl9PtpzXBjx92l4fHvcOUj4P9e0sxCEKTN+/HvS135fYe9
AG8snzy0Srh+1qPMRUbgPlki0JLpkwgmTRI4ZB02LXnb72QZHw8nshH/l8Urr1nI
gqS0rSwrECKjyLePh2o+nBsx8Qd/qzfySXPKcGSjUvL7V8wza3OHkLY0wlOAQ/5p
PaEJoe8+fC6TSJ0sPzWKs4dprZLwlw5fVNlIPK3hls+ATtwf5Wc1kUxfWbIdei8u
GdZuXjt0x5HUJRzn9STXbZc/43PH6VaEwXbxIDOqcnJhtoZRkjcTbTx9xWjBkTBs
aVbktzGhxYGYKsG8WLIBBO5lS4ShwrJNkvcO8D57ZJ7GZcbxfJxoURxOOW8U0BH0
stC3GE7kAvAKKnJljNGOJ9csh0QRTME6UNZT7Utonz48ALanugat9RBuuZxYH4l1
ptRBY1rNEUGUXU+AE7TTtLNzsucoAvZimZk18BWupcni8G72BcGYRlFKUJ5w3ZV1
0NvHekkTutZGkC1bsGEzubxBiCxOFDfH4dDf0bWpBl7dO/0wcI9ydSOigfaztbVy
NSTnnM8O6MVj4lchcvC8KHysMO20gHRYjIqHYC15shkmB/nzm5ZXflwKFh2yVk32
a1sYeb98gl5ZcubkC6AQTLy884KZcX+fCC71TCVvJogZWriKP9EqWHm+PwgtpOtm
krJBchedpmKZ+WbUGX0oaiq+bMXFhnOqnA/WDcCAxeb3+fga82ekudUgds8+ejFu
4NSwnajDHn8pbP7xFwWusE49QB7z2Qq6NxDM9E3G/SGNlJJAEDqywp//SV4cscQl
zXUePPcjaXYCS06mdvi1XzJkhpemuXz6sZzI4kGFmH4mbd+E4FpygRZgXwTGqX6W
sXfVDS025tPRdVTXSQL/WYDgBmen/MCB3zh1kZ/uMV+rwcXxNqJUz3q8isrCOs2P
oa7LbAVbEftceBOk4VjiE7jSed5KwIY73JkNaYCOK6PFCuLf4YqEVyGzaFLhfv6V
AozuzfDoE31z6CkmADjxlALmR0gnhZQBcMsINZm+auKz2VkNYF2movb0J7TUxqgh
enJuasdaq2VIn+pwczj1uaqo5jBAJl3kRiSqR7ATzRy4ElS4Jr4g0+SFJojeQiyJ
ZL1mOSA23mVfvaIXLnkwjEM2mqyBEV0QJxKOEzXAz64SltqW3/u1QMxzOdIHhhkn
/FuCjttMa2CO8oEs2eb4MWPuR1WZ1uYJbTTkCLnkZnsXvVv6TKMBBn1npopx1PsZ
/kim7a9m//OOgcVIPltWdA2eg613oNehqeSNBLpNtc8+tNMkFcjK6isl5MeLV606
RVh9VEvh5XOsO50G5lW2yHsDyMf99VcqQzwWIl6MKuAsK+fCxGGXlyhfgK9rCBBw
FI7HjiD4GnxLkNuTvtifTXxdNy5XJBTFwWmIuOy2uLoRjusoB2cNWIeLVuJihHMm
QsA/Ue5mKo/Gf3HTECHseZTaRasJhkMfc5r4tU+RoHrnsb/imw1ZGFwUcCju612F
9AGUZF3r3YQEyfqELR9G1oe/poCduivExFuT0RQ0XeeqNsaS5Ed4HEJEUDINVaNf
xp101Kw78rSV0YjSM6tutSgVyh95mvcSD1UYfWpAnauorZ4gZhCQPXV5u7E2SSvL
ckDRg5ZWoRWetMZQ2YFmV1n+Lt2dX1GdFUPDoFJLjQkERJgbuKpyYHWETA2FhdEt
O+iq2PwIBA5iBHemnYz6sBS7rPT22JRZDuzEJaF/y3zyEvx4cxZcnKuux3Dki6Oq
7PBFRI4FCG0RMvpZM/3RHRj+0q9YboXLsIS+NkNRZHwx74OHE+r0ulTxFsFrH2G1
5iRxlKOMmw50Gn+O2+bTnV6D3Ozb/JN2cW1ZVBGTsuQ7PSBB5bE2/U+0rCx/vpMc
f+1lOTH9lGbw23EbnlhrPy0vWixykt0Or/vdQqN7q8L89dr/GV7tEML+mYwOLzOR
+8UE3c7Z1UBM8y9aV1/X1ZP/FHErfs53b16CObDGYFTNV2o7i3VokhUp7/LZIXas
Lt0nrMER6gA1pmwYH8CKQphkFFkXxbXGLJGUAVpGkcsyghiivUYymuFfTiwuAJCe
NMkLrEPV5TEN/qyOK3ISqq1EKO0TzUHhBaL5n1JvqEefRqITMbLroIUbyH+7jKxT
bboV+7N0ao/ZS5p1ox/5NVNwdyUFewXzR90VAOgqUzqtUQKqBxyWV+iTjIz9ecGH
31PFVeh5xLs6CvxbhfgGL9Uk6o2MemtDZjzweqBywkvgXbdl0uCS7tshAeyYjXpY
SVZJgX1GScxpwp1KaXitED3PJnmhi0kFTgjyzDm9pQGpFHWcTOi2xFNxobBV9uJK
difXwko95AKJ7dj5OUwlQLGcIFg18/4Yz6sK0xc7YiRrr22j8XQJ8nhpk31przF3
E6KxzLrcWihKCAjGUEIG3T5QrrVnQL0FXH+IuLwJSIPAafCjhxAX09Gq8uEMF8El
DG+Rkk3UPLNp8uLURgqu3dziBAOyeUEsc+WvDC+0LrnuOynizIK+mk35pWgWjeq1
MwikCZTg1y2g4bVyKK1oiMcoRuN/Pb0pCJeb0buVVMVKyr40UKtIjwfRK9Eorsi4
jOcXmsikka0qzihzLxTnkI/nI9jmL36urR5x5ZXTDD9cP0se+2f6HKg5Vw7KRwWr
WJKmR6BCHAH1hNTsq5C6g7Wn9SDMumcQ6Z+pmyRtb5cWw1M5fP4JSsAy1zlEm9IW
DXcbFvOvOCiPs+EA4LOF2MEOyGmbiBrqZ0erxq/J9Y+nRA55IVfuUHFwrzu4XB62
3P2lL0ek8y6o5MpQFpN+BXWG+qXr3dgODpviO900KrMF6Gi/1MLfZFmVFgKEsZJE
jCDtdlLPXG4cp/CDlCOMB3kKCHR7SOD00kko9v8ggny+mZCN3pfGYT9r5KxTPo3p
3/J/LP6bT3m/Hp6hNuzlGiYZhTIFt3kbkoznQBdvAXyvGYel4bt84a3oTcoQBg9w
fAjGCf+9pDh/KwelA9LkM3WLbMUzOf1a+RVZJuxB0CNQNAiWLvMUQxB0ukSvEO9t
GvwQbrFkGVEhu8ifwnhpsjx/+v21StQRnjq9IquP3EaSVVylTkUexodQWzwmYeHf
lsEFf3PKbYDFSuSkR0/ExW63iCvb3MWw0OqM4TM3IcLG60IrpeGuZIXw/9DC3IWB
NfrqHbglGEBcieYIa0QzrZjzMlp9QnNlbN/v/gRhfs5OCRuvdm3np8NZFBxXTBt/
q7KhW7nxIuK+x3RbbDtCNCjKbtsr6KsdG0qXVCEn3O6bq5yHVGlD3St67/drkY1h
bHkoufn3cMShY6yjxu2U+EQ3PRp09Fiq23EbIOCrrHrCqwcYJauDeTxo848Do0OO
dKPowoOtFs1DgDahp1DrhRoHKJ+lsuE60YJNijoWmi/R8g4W/HMcSry5Pe3DwNF5
ba+MV5kAeiTdtPu3kEfMquzYKd9KWvumkilm1w2dVowD34jdx2WamzsaJy6zfpJg
chSDw2U/f7YB0WluI1v1FIXjDf3zYYxc5829x4uc5vDDTLqW++PUuF6mXHgIluDX
NVf5ZGYRVIh9/idZrf3JdMoDBTkV8y71L6Zn4tWYu5u3Ioeg+K0/gfW7TGLqpfO4
I6uPgmkGdN+lEY5IkDsvEgVyIPCNdZJXmAYk0dkhQ0YyqwCzZiQJHcQJMoHh30BO
1Ayr9rB0lDxf5BO3prVmZ7McJKbAKpbIxmdZuI5QCwl9aPoJalAAYok1KckF2wOn
tFjb9k7ortpbqpHPoC3C5TRRGS0474xMvs0IJ/QVit+Y5JEfg6A/iDHLv0H+fTzP
c2pjDe8exSYMsK3MjEPOcBls7swxMt7xn0UxXisbzT5jLvOOkm0Dy114e1LK5Qpm
iPKe5n3MKX2RvnA7x+EHLHH4D4E5nsUpngrS+zpMUN0BcGo6xMfLwREKYwpX74Gc
CpkCtaOHTnEfPx0PQaQk8Iiy6BGpZdmsMuxY1oWiYJMSlLAb7qmNOagDqlCyige+
mknun+/+3JuOfVQaFYcp5ElH9Xwj7T+UYZCHkK82BlJ1BLcTEErwnFrmtl0EIZ0W
AOUo1qlW0pbGRln+p7pSqOV25rNGqKCSRPqWOeY+toepv1xYD32jGgv2wZDzPTy0
wH4567tySYJMnEhhKp197ImjX/ZxPGDm6HhJjnFZvQGjFx82FnYJ+rb8Empes0dj
peLuMaUe16qXv9W3tu7Ip+jm+I2G2L5w7FxNTA6jMv/IyO4qHH5NJHle3TyfV6OO
eiDrVEsJPAXS3t6TFvu+Jk4lVOFM3s2CbHl1Wiiqj3RitAW8hjwn3FzuPGilbwC0
UoqsTk7Ij/Fjom2moU4W8UrKELQoiSqMB2Oksba7uHdxDGa7CiLjbnI/w4r6MPp+
/bsE82SiBU3OxgO+e29EWvkInWKmSGo6ShAeZFsCxJpixce2aYmOn0bSLaFzAWYw
20UZjQLjjcpYeprhiBXB0y/FKB7UffOoi+w+zi00/uELqlh0+r7GjMUOhHkMTclQ
H3krf/DER70wMu5M3+ls+BqrY8+jRA3qwPlGaI4CnggKPHxOXan3wuxK+hPkrPT5
zxWlqaaIYq7gVIrt9Lhq9m7sS9aaXmnPGG/b2IvWVn6p1CWUSibqVv1MF01FKeHI
EsBrDEY7jxWlIeLdDsbvKTM9a0W/aslBrxLkrysr0VYwtR3fQ6EQdoy5yYipvr4p
Gq11LfWItbBo/1/c2CMN4RW6hFcfro3rqvqRO34SbgQ1nvtYtPrha25GMAuIqaJK
9EYj7/5Us/Bme+DDz6HgOcdB15cY5bnp/giuL9gNTchnEHO3rkp4JycjqsYrXvF3
ecUe9Zmf7Uwsh7jNj1+qhQidlkfBnHMJK6g00jpVVjl7hFUYAKUCP2MTXJw18580
OKR8KrkCsjYTB3fGP3+9o25QTab/ZKZ9S/qkVKe+0a9D4VPCUZVbzUwSvIPTksMl
/1R2RRUge1WOjPrjE6TuW0182NpxY9/L3FCsmFkz4imJp42KdilymNoowFLMq5kG
a39wsD0gqFqfb13C3N9lnP0O5m8p/lm+RgcbMqFDrF2hb5jxLXi9MZoNJPB6Nb2i
TDk5ZvlLXQJ2F0zs5GzphT78llrLu3uA002o6xdsfRIVV3q6B7i4rcpRJ5Dd+Ify
ZKelJ6EhHxFHK8R0e/IV5Fu0IVKnfGNh1AozI1dg2kAxb/3GG2lfQfDB0LwQQf7e
mNZ36KQMrMTlU4iMh5CZvnx4AkjQUegIjEbQiunOW40v+j9QZPOjZv98/DWQiuLf
NsCb44eICdkxMzn5Tqh502IwUlvSDSY7LlR2bLNj7j8gADFmYv8p0GJ5KsYQW+Pw
2WTnOFplv7R2XwcNRLOJLF3ok5cs5sbWLP7Og1ZvMM3NFrhk9dggnK31/JFQMrvy
VRnvrGDgI97fY01qxIIzfnSdfVSysCukyQQjN3lmtsqOIgcDd75/s4OJVllQOrzT
1pvC0NG0+the/YFxN7jWIbhVl083KR/AKF3giWE3labCPXVPPuj8BHJ7tUsVmOL2
E+e07Uv38CmZ1WPjSZ/3qrCDBJJh4T0sY4NG5QKBLM5/weifqDDfwUfdYPZSjlE4
0ZqLIi2q9Pwt7TqAZYyR/snkfrC+J5z+iLbiIhfyJm49x9KMdzs/Qrve9ny5JfRn
0hi1Y04EzZdQOE9/JIQCYdWpPaXQgE5P+F4l0r9Otq5pi4neZ//g5ZIrHe1ccuWU
bZx/lGOVgaZNlrxmmc8KlECUk1Emn5R7bs5s4RxMt8HOyXC9X28vJ8DsBbJkRAr0
OOKvcK1QGeND25FRDDAnYQKbqozmZOQoZQpwStVvEL6YG7DuFl7E4gy/QOBfz4cE
JB9Yi2AqHx+WgVw29qJmPNsqG2Hzi/3jrdJV7AlQnqUo1xyEbJmMW+W55leHSE1J
P4vuJGmn/qR1bxPQWBCqw/kqy/8xgf3jfKiiuBQWDSle53mu2gKl2VyS7a5590HF
q0NtUIGiaReOBxZAFUHqyOc/lpcbSNWjOV2U1mAr3mGRwuiCFRgQk0TC3/d0gsAN
yZIl0EMinXVt1k0Jil8WBgV+pl4mZKyoPsJH4O/GL+FyQW6+RuBcUOZGSxSdAgn3
0xSa5lunhxyGvar6rSxPIv1eWsw5sQxdq6e+hlgUk6i20djrGxMHHRwUAdF3Mx8Q
QxuF/tk3H22CHUiqk2bgsB/n66tfG8bYuQGmUQpF6fOdMqBBQx41cjgvdZozswIK
53b+8ZrWtH6RW1jdtUqC5NEj3TZWP9mQ/IkhT0EtIgx9ucTSpSnB1/lHbpAaSfgy
cnm46uXyei/UkKfB8KFmZs/cmYl3Hq3Py9R7Xdo5jmxml3xmc02mcNzuOIEXogCu
LLsYS1E0L4FxPQLD+EN6LZYFtJ1DQAH1Xo9xisG+v3kZnD6J2rgFUnMU8yK7W3jw
YBRJdBeqMCCCqIaxEI7XWay+TZdAz/YAdTnMiGEq1MIzxxEmsGzRJrawvwA4HHQ6
LRogKKtlNNAweYYemUvGDk5/PuNQoF6G7T3wGH3JsNsBFe3CUglWDB6P93QJ6KR7
OKNAFC8yDqsybpU0kgIaSmZERMvQcnecEQmrRQ88XygRg+YkH++IIP69SlzErj6a
/Fmn5tRZPPM2mYocr/o5zJ2WcyGTwzqFNOM+3NKmI5zUadok9DR6saAN04yPpKFy
++XUDu5Jj4SrB331nYRMcyG3cKAUOrlstSSkiXfTrjfblZcmRjhgaPzFNnEE6CfL
Xu+IAcOICk2WBQzBCvhpW4G+b2SdO5AInx/dncOzXqiK3r1mW+w3VGUpNyxfbKk3
M/8tmgG8BkDTcWWyqbIJ6J+dUrZtcpVjJqikL64pHyfoycab8Nlx5/LZCcqbTN1p
HCHpUHDWW9ZFryNWFk8S/3KVm1M7tML81ZxLedIyrNFVQTDfdm/wyOgvFspdQr8h
huePtqTGomZrvZRK/I5sWv1tLzGEe8hEdlE5vC9vkjypdJgEjFpa6HIBbfr0nndq
KiGhIlBawBsImxwyYWhedW+QJZXQb2Cfj4+MvbtrLYmvUKvTuZr+Y9kCnhzbdGLs
6U+344DxL9nf+E32VOFwoRXkz1uvRnQoB7PlzFMf/XXxpYj1z5zsglunr0jf+dTq
iSqlFpaNoD1nKFOs99/t6Y1Vrz7SZOGm5eDrKQsXUWIRMafxoCtX6lo5hLml5Kk7
Px4/ZmbZF+1j9XE+17oWu5UGplGq/YrcZDo9MQrivOeGraDDFJWAiCHKuKm0V1Iz
0zQXI4ST8WiCe4M8G+u52OaqLeXJKZkEP12fZCBYzi3cfkM+5My1uatE+wy4sCCy
VPJGHmxOTn08V4gXQi8l3piyRIdl1jt7Rl7IguyuCOGXKn6Ykpngwof/Wqt7DQwJ
riZY4LDU7mh79ZKnr6L8090u3TQG/AoiMxymfx6EonsUuOwkUpKTDv0bh1OUpzzG
DwUmPs0Y4iM/xWnvw9SJvqtk8/L9vrrsOS+DuE4cREWIq5+YB6zJ1YUvw7Ib4hDT
FKbTnH/R3cC3Etp0WNpVBtY0w8dnXRH5Os3dfU2Jb1vrWI+wlj8HeZhyrhNJ5sr3
YselegszFw/SOEGnv2Eh5MjTXZgBGkZ0PlRNb3bNLiFvOrWZj572NFWbBz1JFsFp
ohwvAk6W63t3s8sNTmyJAPunxy1p7ogSQ3kvnvS0Ewcq0edWfzpAnzqH1j394dcx
pENx1DQ0DAr2iPFZvRHkRhFhi5EGc0HV/O1LyYX+RH5HedvTSX7nJmfFBJ6THaLx
ICUpjmsOw6/BsDBk8ZaHmYxwFGLpCxZBDpxwACBWfyymgASwSMooocIOu8Cps4sD
YMjQSSKgfhQffZhPnK1Bw21UiIy/QUQSh/d+wovQ4xXzjGK8EJwPbyexfts4KCDW
TsoafwO3jHqHsETeTcDy8B4d26CJsRqnXtCHRufI2fVOmltAmjRrlrpLaXGpmPjU
Nly8O+ai5P4wv6gNffZ5X2ssj12JHLgYfiNhyueJTlF7yiNSY2zM7jvlIkxeQwcR
Jr2elgviDBSvhKMuKmv5YAJdQtpGKLGdPlx61rDBDrIxiSAIjOLezwNnxOqx3agw
udEa10dF5SqfFPXMnJSZNlp1GOAwfhKWfmzqjK6GCeg93cohAoz3hjRr+dmyuql7
1Ahmc/9Ux+ei7E5xebBAa/dYJoZkOmBxTe6y0OLdY/6G+uprh5vGooRGIza33+JU
MxghDOtAyD+b+eBxIHefvva53/4/tIi0m2oPvDqCSWZOG8DvuBL08fTNTDPnRU+G
k3ynpn83P4qqfsglyDNCZwCHQQuNq3wMl8y+kjTSr5y6wVvE1Ao5ZOoonjjXZ+zz
d1Rzo5+8jgqJK3nBPkH3pLKyOMidHM+2OFjFUnzfwdC7adCRK8Xx7a83+fMwvFtA
9bqsNUFJB/e+DdXuowjio0Z9mC3Are/nGpkITvMxpBXRLnkV0wbyayheSli1Z3kj
UJOZRhTI1ck60E0TfH0+EtGoWuVoFVbTPWRl4+FMUAFNQCkOx8dwUhWDQw/YneAy
8+r4bq4lSQ0KJtwj2TvYvd5mPzNOwFKOPd5c+YDvSjofhn1KLFAlKMnbqU3A6TCp
XXxrWXKd5OArMa/w39x6TWj5NHx0R3KaaZ3FZiYCUj+aCz0opBtxNyXHoThdxo8A
ZA8lDfkB3B/V4Eb4rjQJmfqfI1Vgxq56pdHTFI2NYcBDDwiaUfzT5QxaBw7BnhiS
PbEhWuGRrSB+mzlwbCKRTw8H+E6+ZFNQZ+0kZbcbW200CfrOmn+el4vArmjZJyXK
n+OCYh/UIa/BmlhzwtJrc+jDHm15u0eLdr8hBXzS22aY2FdEFiLAp/4oQa6U5TjJ
ChLRDAumPdyovuJ/v/TUrm2llrfJs7jGh5QYxCoAjZdIR9fHH6rKJ/OGUVhdI10n
OWp+fv60hbe+eAYfKuoxZVZCF+ketoMl3M4vBstkqx+er2hxmkF7b8myZYIv+lBx
guPMbAZp6gjUhd6dbqwGu+cUeyaSHfnp4P7PCbX7b3JxrA5C7fbqesbFp6AyHgVv
iNlaFID2GanOs9xfBHfARKk/BHkDw2zuJEznkepY5z4AqC8vomos0R5P1C1QlXTY
2l1ueKSOJKxz69WgW+etK592lxEGN+9lUMaEHxoU+pSa9ysNynhCCY8KD/uwSSaR
AY/9waM1ZuxUIZ0O0pn66LtPht0sg6rz76CD9LSsY2JnjRviNoujDvKKJSAY4Mal
X4BotyIAOMtTXSiwsHlqHXbfXpWk6A2AvWUbV26K5CIKel3QjI6Qwh0BjkIibnti
2mFU37khc7FL1WlE/ZKmN/ZxaIsZojyedrQAUu4e6M6FDf+vYEi01GJcPTAIyAHR
5ZAzshRcmzqxCno5p+53wuzRpNC/aowqXaz6+YsQ3Qsvook1cVPoslL5TMOCGzfA
+KjbshiTxH6ZN0L+NgAwczHWqM1fj9ZtHEfeQSw1e0z13yKkqCQn7Uwo1v7bELid
Z6kGD+N2W1gA7b2yPQUeQV1ahc3ujTb9hhRskMh/T4bhQyiPMEge6Jip49aBmDwo
xJ00pWD2VgfSr3sCe5Qfl81fGZKMEq3u+dDQOiAOwklb8BczTURugnB1mPld1mSB
2ip1Dae3scim/0wfRmYZZzJqMDiXcPEtNCeWjYvfc5HPZ+SBFT2Ple6GfOsmVAza
30F+oT2ZIAEzleRzuWHlgNzrgrJ4X3XxIg9HYaRFRU4qXDbEn63uYOQn4tdQOjsZ
nMZmwCaqunxbCO/QX3AQGOFirkQ5MvCobInfWkD/w9aTRPqs1aaoZ+RtTH0CHurz
6WgCKHz9wqMziOohezp2rYrbh8THr3MfXS5nrwRhqJJrTpD2zyYdhWA17dtqKoCI
0Cm7Padr7FpuM6Hrog9ori1STUDgySx9nkzeMUyMNtsUJuuDYBAT63EneTqxKYto
aqTwfNBCJcicHd31C5yVoSavvViroePtHlfqUGp+4aKJr1FmAHkgRokqX5VMA+7m
NVrlD3JlwAs6M8diOHS1eOhiBvujLVGLuUR9RKByS0hWA9yb4FMMJsoszVxrxbin
lZ21+03R6s42gDAa/Ed7LdLI5Nfbc+d57TljTZKrEGZDBUylmU3vzD3f4Aywzyln
lp9My81SGuHJ5ShNqLs1Lwx+UtEab+T768xsLd6MNoOlmH4x8aFQDLhcmx7Ay3Yp
INJykpZFvyl8AorkcUUGwyQ6mZkakv12TS2qIM8YIbmCuqR78kBSIDDTeOhNT7pB
yar6mDRmhnbI22NsPJkdsYO5z3cZh43iY31XZywmVHCoapqXsBY+gC5DV7+QXQkg
etPOsNd11ArLopkUn15RmHmZUJaPo0NwAq73cOP5Npmnly+S5uiej41QQsQE65At
hWclcGOXXk8CpPgDu0i+3k7jtWRJ6HD+pHDtet2YD+EBya+MeBmUhaCHQdqnkr+n
yhOtZrozy4q2giXXeRrNbjNofefMIMtk9VFL89kBNnnOMUhKBAkNoH4TaxV+Rp+o
yeTntxlSdyKlZJeAIwSoYN1fUtw7epMcyaHA3sDB31oclZ3Puvo/mz9kGNQ2PwGY
c6mbX5lWImCt08TVeYYGj0g0gQMCmLPwYjJbbf1KOJAW4yM0CwJKdiQkDdWIKYFH
0g+RhtFJki6DSSJ8aiY6dVKz5oisj48ZDNSvPC/ZVgZ2iphfDVY96YNs55mr9hqP
lgWqzoPe91ULBIGalPqa8n7buX0s3J3ALiUqncZm7hIZNoxBSIaQVA0zTOa2+8FY
p951q/fcXxN+oVzXATfReSkAov25IETzkIDg50IO+GscVA7BQTrFis3KgSoqBMay
anavStCs7mWIHOtC05uSn9x9oXNgKOgSxTxjVaioafIzSZ9MYhIWDS2y/47JtHj9
NzYfV7X50qYYPrOAD47a4TwKhEgZjZRVRE/3aWbx8gTVBDJKlJdmFtb2byEe0D3A
GKK/kWy3FZNEYRS0gMOSQ9ncW81UsvzWhWfZcgg9O1ILuHX03J/lHHrRuZtkjA9R
xP0B6TFDmZFXGxX0M0y1RYjLTsDEbBsHcaqR/5Pi8qp7RP4xoAUCzMLvbM++8Uk1
SecnToRMPRCGN+0BbgwgoDJfhg0DNAq+2I5xA5I/gmN7o3t9ABbYKg0aacseJ20a
R7MDtnstIrslUQzMnmGewu5tuB4QeQ1Wvc6yUYMQ8QZK8ueyZ6o+mCqp2fjs/jTr
bCYztsDgTeBgKwBP54kfIcLd2Odko7z/VmECbA6YdY/JsSjVPm0ux1GCve8TxWvy
F/lscQQTDJm56Qj54C7mSKK1u3FONtBNCKu1aWsCiBbmiMVNiW2mFmGMBO+V43LA
7eyPjFjPVIAL71f7r/UWDc7EEMyBPuasQ5I5Z20pFxighpC4rye8aRsv5uujebJx
RYM+NMlVoPEa4vecT1/pR4hBbkmYBWteoiD+PpYamt/3Tutb9J75TP52II0X3YNS
SZoVyRRwSmVtg7YXiQOysmGrFF2eHnpLRyytVr5agFDcc+YX+4eKLxL9HrE7m3HT
LCPel96+nlktj0yAwqKL2HyzH1yWfy0hh6bDiXgdDT9Sg/LPIM1fgHylI7uTgHZ3
RLJPieNiatcEngd2j5NWO3yf/XkWAgo5PJIqDJG5d/v/86gUtQAYhW2aCsEF1M4I
Je2hJdss5z/8ofFKZ7uMRJ4cE6iOESEJQ4u7niW+sHtFZnRlSuTCpJFg9rVAI/QS
9ah4UtOd/XJq5kT84pJiZypXdgMvVH4kVRwHmlGTia4kUQXM5aVwoPhlGCc9IoQR
qRVvyA/Q3JokXMvuQE45jzcP3qBJh2lzZLnnLW31KXSSLNfian3gvYZXAazsmfXc
XfEDN4VXOWg7ax3TfgdxZlpacCirWr4FaZ5nHocIjEZZY26K8p1rsbr8GjwwtLNX
oSqsex25OBEju4AoQU+QTQVh9yOVvFHb41zV0/BVt9u7jwEdmW2AwjqNXaMxo5Dp
Eu/pCFfe3HJlwgBd/Qc2iV4Rug6NRwsPwfnsysEPn6gxqjq8AEnDgbffyCaAvAkO
2CFrW1zk2r6mBTn+kMTS/3Snlr65FOFEyv0C7WIVagIniOVqFFAC3i5a+GEcUPlL
FFPPIcZT5ZXVWTLsFoOfU/eHeDOIEithp6RtmpU+KxScHlswl4WsQpHNZUwSwrBL
ox8uDMp+/PppsjumnMeruT/fvZcQ2pUE8kgBchi4qdd07S8zwg+iBHXLu5sLdejw
gMzykfq5y0zHt5Oh9EawM64adNIw0d64AdMykR+w4D+z/2QXR/+9jrGcbWFmwByx
tXBlVOo5HNxwcLRZZLI8ZeDJkvhGX1oFuHK8EuLDqKsMcnZNdwHgjsmYZcx2NuXD
5yMZBpMg7ao9DlYmwumBteVIEMEe2+eJLCX/on9Ap69kDtRqyrYv9xw5dShUCzQV
W1mdHXcRk0V+40CguVnto50OL2o1iPFcCXihmDSKLq1Xrjb4bptSWYOtbGIeogF5
33vuiS4zxX8f1RlqxoOxF9X5nWtrnPxJIssbDPHAtjb4u3CqJIoR+sCiOn1rCRi8
HdzSmZHhy+I0BqOLLKq5u2JtP4vx1c3v2mm3q63FfiY1oxgdDEsotLinJL3a5bsd
gaZSUDCP0JoA3itxcOq6NwQT3FDhz1wiYdGIsppsI0/X+8IVcdXenmaq81MvZb2a
f41FmQZaXgtTQ/tWbcK5Tr06hKfGyySucvVYA5uLD3OXf9rpdnSIlzpy+kPNkc8b
YYRF/UG8Ue7Yxu1yz+a5lXVRY37fk84dmPO91T+pd0784ct2+q/RbdLaPsNfsnv+
8fm2uaotKushRq1wblryewZMluNs5zZMQDo6ZoFWt6eKNpg968UUOBWZUtZIaWxC
4vmebRso+9ncmZc6Ot3koLAugavrDBPKWNmyaMDEuwnbZtbcRHg2qTLfq2auTMwT
b02pG6l1SnddQahykZNGNlZg12v63l2ujc7CH1pvf+t1QpYeo8d9ozS04Z80sAKY
vuSJqZ2gzcFX2mhWZpI2Ftcmvcf78/NhBkLtH+dJAD8NW28PraZOU2VU5pJ5kEEV
QYuPLJzAVvVOPV1dk13rGSAIKUuPYDMj+l+jCl1z/IkplE/XazbGjUstrTxvNMMU
4nKOSMkBm8ELauqWCpoCWRr1b24pkbgllyKGf317uehEiymCTDMPX3tQIBXG3/jn
4vH5eXTvHZ3a4ggldj4hNvSA2Z7YVj3iPzbpgcaT+ZOiqPNSQp+/q0lnCefex7g2
eajb7ZhiVCX8C+Y3fWucT/buPTdSl23JCrXtMxcxTQ77oT+4XJ1WVzt2+T5ufvVX
gJrB4pFaYGWTU3UNJuxg/RQ0Y1PGciQHG20OKWK4ZXCAdqcpTBiAhN6lvPo3I4vI
Sl5uXPdGBXbcU1kJs4Swzfrw+dN6GkgZ6Xt/59atsHL8NDb5EbfhaSvkbP0Ss0jL
GI5+J/eW9evg4Dc7GU+1UjSgdftTmRCjoF9CE+jOugkk31pYBiupHkU7bTHiB3xa
B/Y4E+JfYfb8NQRaBxdo524a9DL+q8Nw8N8+aFSgPGImT9iXqusManKLpxWNeLJG
CFpLjzWcmNDSS4CUVjSSfn/vT9oM4vPylMPXQqZCRyAUqaqS7jM6xaLjUXH6PU/o
b0k/CFsIYkyG6m3w1eYadDo68I+5oonSdTgV/Z7e6uTMFX3JEWzL9pu9pgxz1n5l
7DiT2JgryknOIBZV3YGgqjlZKT2VKh0tZXVKCjCBU/KHtKbeMcYF5D+QzrLxc0/V
obzaZiiR/VHII4kCcdcriisrc8VQ+me+VYjfgoge/N2gbX6S/3KMkvwU1YbhYaIg
+jXjLMy0eNL0zZpEeLdQElRZYyT7povHUiBGUIHPtjlOEbmgNQ95Sppl0Y1/oSL+
a92pzbXI3XYG9A6DGtR/q+3fZiksjijePZ5gd8AnVO/X71QmnVavig3nulV4+VAU
e6Fj2oTp3VQX6W2dRkIP8sIB5ml8N27csvolVXYfAoJVrfxsXGPSadIIfwldNkhX
SM6PQj7O9DKfKyw65ohWZ2wtHxgOmEbnQdsEtIWvoGRSg9YZYAEWvKq6dAYJXJUV
AEjTkGP3ob41XdCjH1+KW4NYhhFgmvqpRjuhCL1BaiHqnoDo+A5YcnU18XyBzUpO
/8TsaE02ir6vDoThpJJpBU+jMWqhjQVtVbcU9yg2SmoH8Oi3gwnCOOvChxf+84BI
RnngO47PxNtWNXvtf6953M4AoU89QAKzRYh7N+GwgDBnt2LF6SBJT5Q6sAwse1/j
Eove3gDmMSBiAQJhTU/FPOvIZU+8uNNMI6aQRIC2Re61LlFk57wpuxyxtBafoZXy
TVDUHjIW6RDCSjwFToonJYVzgktMwzzNrpDxk9XytFISf6ulUgfuxAqiwx9m9YfO
fP6FpCPdfcNP34QAdlw8kUgfBy6y4TGgWIf7dCR9OxMh3bkX4nqo2uZacRd8L5IS
2lALXJFf8pZBDilslSdqnx9j6D3zMgj2Wo9RMWs2kKoXw/rvqu41wppfTA4TZw8p
B5pQLF1DYwriRE6Ho1T06Ahvl4Z4kA5EgnhHrzdlG1bgZdV/7jrrVZFprmBptlCb
INpNJ7EW/p3IIsh5lt0jcq2F1ITp8PsAx7v3Z+ETjbT317agIsxvOaOz0jB7MjjW
Ux5RuC83tqAKQV508ee/pu/gGpocs6tPQZ/I+zR+1chVabKiLHMa1xzXDMMGWETM
Rryd/eN8XmG+GPaTkoaTnJLejgUIKzFhXieOtJM567aQ3PjhJVIH5EwOIj1VNd+e
rxSkq48q35HpeeWKfSefs4S/ws7rM1zWIhzQvfBxP2jXNDq6YD2kT+32kDVNuX2o
yjCadlQZTXvoj4nf6gMnUZ1Vu/KJoCdHIp99eoBz+9s/Gh6CD/8pxkwmOwAystRw
KDdvlOTfNzVI7Bf74ddIBSvUqwGWpo2OvG1Bg3zEI2q508cqm2hkeRO7c+Lns4GX
Z1CWMJ2V3vRjI2mr5hLwbgF7Ol1+5kXV7wIHM30RHmWKrIU0w8N2+7uuJ+hkBZjp
C5llw2IJLoshLovPV5LV87pm0sN8np571Acdz2F2iNQUmryhTBZPooZ5692EtX3+
c8kAfClKF1Xqt2GWb1MCsJMBCfStrGFv5+NdSK5zTCDni5bGa5ykIlnWVH3b1ThO
MCo7KirZQyif4Pxunf1knTsmF6Ij6CtkPH/WUoByKLlO91LsxK6ECxViLggGnMwp
2yhMnvVvaVHk//wfjndab5xgc9jgI/6AV9EcRR99HlvY1WWvCcQIDLyzICweQIE8
9RwI9lJcQNLf7iOrCsyPHols+x54jGPHrRpXAYaGN86TgXDpJLgMVsMS2MCQ7Nyp
DHHcDxxDW3LmMbTlXL1Fc1ea4XkThfW09lqeg+CFmWoMR+cn75ob1lOXwAb0ZOiS
Y7cyjt+xAT+2HbmMMtTrUqYUr2DB0JAKka+pSy7ZcNtmZIIPVMUDXx9XMLyuxUbT
jutuxycPAbsj0jZee10CE1UYmXQ8y7FAVJYmSKKQvnYbvfr44ELTO85/BT3L82I9
WKE0FsXqUkppe7RBGnT3CioUztqkLQfw+A0OMy+iCEAF8EYHZ/uIYzFa72wEOJXP
3EjleGm29D2Ss/XOGD3qqHdmXojbwYALvuU4pcRXl3fYT/8rO2B4pztdrq25ikhO
HMddB1d2+BanUpH0C8Q8Q08uHN4VyyBT0Wb+Jri4DHEFgZZ3vUl6SWLwRRbTGJWS
zMmfcZ/COny/6lQloVTuGFs5sR6rtBCwLkAAJfEL0Akx4pOwQhj8ERPswB3nPBZK
BN1bUVOZHU3xU3hgoVDcQL22E8Sk4jBtNgar3aSURDLyK72kFeaagggeIheYsNXs
XGU3+qE1W3UnSZ4KNmkShTLflcllSdV7q7tuCHLQFqAdkndAOvLF20C28cELmO3m
l8Y33d7WBaR9pc9Q7nWyAXyOo00CYiso0AysKhB17iqrD+pZCrcYm/r1GIDpD0uQ
7PXSX0dWnvAsbVEAihpvaWOTsYbm89IFzNyepR4/OxkIc0/EwDv/I6FELQV8EF6m
y3OnXzeaGEYcbqgOz57B/T5AeBxqet7eoaC7T80SMvMh6xPlM3Qf6hkphHlxXAbA
12ogjPWKxyd36wcGmADsQps44WRpvybhPvagLFrz/717yLgpdPWXcc8fc6uhmx7a
+NfPs2cONTn2n54Prm5wyr/xCALUV03ZjSwUWehx+2LFIgWw15sgqmOGL6cfwHAW
OtqBQYLUrIyHsnfwMrvU9Ow4niEQ9T/vjsLXLDbkbYczpUu2Oo+E6t1X42x7Xxux
VYvA2siZLUmcQaciBitpGNBOVBs6e9N28M4PFaU+6gmmX6IaxHSiR8PoFvDq4pPz
GQ4RS1k/KHNutb32D9j+ENzk8rNYajaYEGdMbk1639/srKkmNBKAzGiyOxgA5oYz
rnAs2HWhse0pEExDRdq060a5p6bVhBU1/hnS1BjCSrNy0Llw4flju/dahVQFhz8J
qfGtqQqZbdD8wuEsAR/f8JU9402baqFtAj2Hit3jBA61gFAn+0YA2ByZvdzTA1jc
xP9Ros9XH/nj9LiA2fDlt+fRcf+y2YNa9GIIbhXubFp+6zW2/JI7Md3EIBZmwuQY
FCJMhy7MjCaBCZ6iMlcZKuhR2i5kZnNcimKM30iVf6OTXV5j3TYTWQICnIYJEpm3
qTT/xdVL7WUlsGGRJWUh2HNu2lt264Fs3hbGXLIAFSEskgSNdL8NjAhyBp2UD1MD
kTDZ79ekJgxjmpy0lYPXzjnqzXBXzeGUelPtpEdJq2IbIKwrb7g0ZQTp4+DfwqP/
ry554r714WTX4We4GmgE11dTZl0c3gDpsnZv3hXSnT4OZsNZDTX9VUtMbdf+FFkN
WSCE6J5LT20R7VRDbxiL4cHWItluZEPPgUkKpd0OIWZPfKOR/s1pm33Tm1ggkTe9
MGxpflqpo4hpjU+mWCWbchQgCeRalmUDZp17f4cJPOQXvDEnIqOTJelHgkOMTwLy
VvU5sjx6ZTy23+F2qH/Ci2kCvZB5OpkVM0lCRSLbBZbH1Nrm92VgboIcwtQZxTdY
R6VzV2Igqbgap3vdPU56DXvbTzddyLi7OBvFKDSe0kMgGmJsbVhmA5tR0QLU/u2Y
EuxMvAegGDcPYbX5l9mjPHjppwuyT0YHSmV6Lkz5Xo49Y9vIfCkZE0ZkZlkF8mMf
S2mmt+sLtJFuJJXshh/+WC6ojqSaMmbGXl0+b2Nlgrp96wA01ZCg7cTrUyOZXyAK
QQuf1Dd5Lm408lO2Pe0gJQ64UYv/fFsSvnKZka7AfmzrErVXTU6e5t7oNFEVtoXJ
rUitgAzLk0f0isc4nmalVD0z1do7nk0vxtHau9W6Z9mBs5/iFriH/uQ5nQj2NgVn
03h/j5wOqSWWg73nLgTcduzIGhJripUyJpARY8WdYZbwOwDScFdmJVHHrLVxHUqs
IlFW/A+DXjldJSj/D27Cq4YPpaZkMntKUm8PA8LIlGcwpjhoAFHBQTStP8z98kFm
qlJvieEEUsJVBKHzrdedCSBO4aqQc+aCzNWMj3DdxTnNLs5VYxbnYGn3cfTw9JDT
Za86DDQFh/Jw827O1y3pEegx5haD2eNmJvwjNVAr3gic6HOeF4WqXvEdFD9hzrid
ZfcPP0wxGyPcHJttG4gyRNmc922EMDqrzdF363tE8s4OdG1mYmpN3Ib6WdQEAnaO
PfL2ki1rUrEX419crtLNpxgHpY0zHNwtuoPHFHvlvJVaegzimndu9TY8pBwuGcW9
oRm/KQZNI6l/9b4WWmlcXyZP61wDsKCiQVrCEn27kZ4vKFTv7NWu699YzCb2n5yI
BjTmnvg237+pKktyu2RjDnrSrti9Em43ExyDdakKMwEGixUmOcGnrAfnhCCVnpd5
X2UqjdE7K9bQIVgBqhaQxU7msJyptQUisX5e7dK9AhEsl3quxgI6c/AIrfiod7t5
8643S3Hvo8w5vTLpSLN/hYlLapGYgtYe4Bxkx+7fyOLF7y5faLErXHMMjPnL0WON
HvxxyB847lloidcqa6VroNQ93PGrNx+tNWIuN/kHcDIOHUqKlLYmap9VxZq3a0Tu
wuxCBhZSIxvMn0Fb3uBH1OD7JhC+KQ4eajAKGL6H915c/aYyy9P+l4BszLN7IQOO
k6PfY/7ndpHBrdagfGfVW/qrOqgcn3s4RpQecUCcPMSYstTiGAXAk1OnZNwl69UY
rAd5rH3P7qbC0zXRoKwc6JHgodHB0QaEwiQO4GG42wVoo62fGgd7LnbBO6Hd8g2r
VEBlPLg7GqRprCKWQRzGvalRzGtDP2fAnIouFiw3jt8ajpoZVo1ylMZ+cfuo5BQg
BtP26oU2WHwi/V7WBHgpA2rwE0RflYTn2z32Dc1dwqXgZRCvb8cgS2OWF1pP7svi
gZOezIJ2i1RXK2IAFYVK5eKIx+aB0Be2CfbE+DfrmIRjB+mEyaVLwOTGdU6Z3xNO
pLqFqcgN8W5p5hzydyVSXg8W0UjmV9Sb5Rm5NH9xH+JPgG6/1EqdRHX/JxE4VP38
mynu16LXYdZyt9+LQScLYNwQbby1jY/C+pPHb30f5f0sIfbt8bgEGnExFmFxbGIU
NDF+GXB47kaqOTqvisQ4TcsHtK0aI95lgAeItQMzKOrFDLszUPBi18iSYD3e2JEX
SK0zK5s+kVwQVOIa+APhnLGJlScCDzSJgPta56252m4rOn8RTEP38TemrwMO53ou
TstmHv3w+0mMTXdmANDcPt8L79QbsFDdfN/brPvvvlBnkZxyKAcSbRxS55Ai59M7
kwRRfvpWSQBI+Jb1a8pYFvM3/xbTS7M1dRVJfw/jVbPKkUBzsCCUYUNXn4DYCxis
cxZ0AdgRQJt+j8C8BZHi3Mk1o7G31z45H87UO2LrNwlI+GiIUtnsdZDV0Hylw/bq
DbK3KjHQv0cH9YMJWlgg9UOIoc5aSqIlPjTyHbCYoHfhHCCeioMuWyOeLZ10slTO
CmEyF8/rvpa2gsgDKpm8Zi/VGmXCbg73IKgwhvWNchmLDXO1CsJFgT2tsdAaFzjd
FMxGFHBDybMzYMnkaFm9YFI7OdslhEg4mrGSvkHkXoINfjXZYEJhqMJ0jVuhCoBO
b+vD3FlfMOOGZdhf74WyR+wFGg1e8gcFj8GOXJi2gDn5iTIe1uZBoSldwjbwDYJT
kMNc6/GeUYUOQGoV5A4uT9WF2dpeNfX0Ogh0yfzA1aw3gqyP/o8nWk545nwROulk
ZvNI1rLhik+1Mw0yyiWud8bRULeGjwXip+ReRsGt3Moed4aeunNejRWRnQuWVzRg
WoIaIVtFYhTl3IECV25DoigpKVziXg8W4R18Rz3T2vGNLUBXKmj4yNOJN+4w7IuH
fa99fLoiJIW4U0dqU2ucdVBjDwb9klV3X1gY+a+lSNVW6vTPs2yHi3MVHlPU7Lhk
P2+CqiadvMjycT5h641L2UY8p+a0IfodZy3/UBizh7mSluPnYt4l8jv2IhrAVRWj
F2SSb1wkhO3D5cdbBJhWGFPlDD6IYSrwiLHCAyTTwW4PbOqpCWY/4T4RtSdTB+Fe
iaspJMj32E+ExRmOX1L60l+RgraRrabvVZhn+Bfy6KjHfQkU2RiZA8kGOrwxADVT
DCg9ePqI3mABx7G8YJFh751UMQ8es1XSn8cOJEsmbp40UAUMoDuknOeyT4WvAGc2
X8KDDyryboW80y0O72BNPWQfTsvyFdDMG8Uwc3/AzUtjYwM1tGoVbv1AVx5T5pPm
qk4+MFNctK08oTgATsa+PtPOuY7Gm2+z3HnsdsbIcH6yVz4AqMeRvgyGLuzzhAFv
Jy5QRPnowAf7arYtHSLU2CDdssMtwm32oUxXsRVafaqQZEX84XKoaCwm/btcfo74
Ni4wquGJnNthL0vEzBGc/6Ib1hTpKl+oEe+JXpP+WnXKt3xWyHFde7VNfI5vcEwg
gUm/vohKTMEAX/rRm4NNfs2Tc7LNP3mXFtK7THBcI9A7eNvwQGdG1D8LbkceXx0J
4LDmZf87eOEB6Ve5+eClEs755wvchmCWjHkSI03Pz099y3CLvKkN2Z1dKpuvJI9z
ogZK4qa/leqfQq2Ez+cNHfAPppGIYd5/0Funf5cL1QDzVsl5AxVPgd00YG2xVxBD
znI/g9A8r4uh9+40LcVNkzv37zPKzTjlqkFtxU6RTwewhEAr3heVVdAVrvAtWeFO
AxGUPlcrrL+OX/sfN71dvnNN+S0iOY+Xp65wrJDmExNa2bBNsuV9VvXyfuJx3C91
GEcGvP77/zzkmyYrIfb6cGvvb2AtpytGk+U+FS3L/B5qzhmOYRe+1AsQ3DSrXBZp
6ZHzUq0DKvWS5cXyp9UuMpfV+GdCn/lflVHXsq49KFeEDWs/6K1uSFK2X3FssrKq
XrYjUmTSbfDdUptvf5F4BIW0GxtumShKseZ0taxFC5NHuBE6+gYuxMu+vk5kP/hx
yatgoi+/ObQ8mvSzSDh5o5VJbX0EmBntsAx+qQp/9XxPOVOGJZGQ6qXglBAxi3YD
7VTh/c3CL817pzshfdfTL5cfmAAs3LiRRK9szgBezEZ13zJ/cQ6yu/8GwiT/TZ1c
EGeq8e1O4jxqgSJWxCY308//xEBVYYMDhPp+0U/TO2T4Bj6C83VCRcBJFwFy7hyR
qRYZ8JkxmgbZAkuoCMF5eaK8EQwfzthauNnyg1Za35VrDRAJ6csntRBBW8RjfLcj
vaQ0ZCjmGqRIeHYSfM3lTqe26B9voAJ8rDzPheOLFWzZvaYRSEijC4wQ39BVct+8
dzbGaJkOKGGSbipX4V08tB2svskMgtw+nNPlNlVgEXWstROF3mjKsXPt+LwiDwGS
0Zba0e5ZyA0TEDen8N0MaRZdrFk1Jtup+TvTji+bCF21EGrrEth+Fc7Alm+LuVMS
96X4ZwQuFkTFlGTmNpvgA+2u2Igelm0MvSVbT7jmKXJHifUwFs3f2BW5U05GT+qF
lb7XoWfN/hQD0nfRsr5ioxJ3g9i6xCFjpGJJBwbN/1P/DxA9oLgcV4dosUsZLhVv
ynQMOxESUf4PYLMQNkASi9uCt0pJMWj6zfoSpyaYM12jOB33lK3NDfjgjVv+Uix8
otymUM29thDiIK6whJ3XSJP5zB/hfvSNxMMBNyyA3PQTTFGdcw+ZnrStiRl7XC1o
9tF/m2H7XOlJs5Bu3XzsJLAsVIPXqSDalU/KWXgHqZZKmWoltbEvmOhJOpfrl6vA
BtG6HzmvqR88I2aedeivc6jYzI/p45hsIHg2X0rznOOn8Dj34UV9rwxhQpRH6BL0
qsBzx7Azxr3W3SqrU+muAEvhXO8xq/OhM8WurlbTn4D25jZULRRUY3BkBDOHLIji
O+/31jwiPIc87ATRamCmkqz3MZLPC7+I2p0AlvgEYlzbhLG9wb/q4s6bS2B4o+3+
HQn4IR2sjoqnnn0uW4DwVmSKhuBOCM/0U5UKD2/ZJQ3TypyNXBix5/9tqWoawbNJ
QRYJvVftWPIEMMmTsS0L4a6NxeGuW78gOqFLmhwVJm5oQWT8k9yTC9R5Bi8sp2Tp
EOIrWyb+baRuh5Q91KkCddzHp7IBXLBkTjwHkcQ8iIYZ/sS2n1Y4uAXXkD8N29zG
UAECFdGjAnPW9DPog9PL6Velxl9gFB7SxvZny5UsWiXZ7vpjMDhbbmSjOqZnGe5J
FPFx0JYXhQ2DjyHjelFUPW4YJfhksnVAP27sZA0ktIvqMp5w4BTl+e/+GsLcz7c4
qzhjf36BdNeKNhucoj0V2yKhkjEr94QwIUFemz/C1KG2xkXH9/Mh46KMxY9FVoMP
T+1+G3cY/NU49pzkJZV5ZzqbKQZdcrgieA4l5foie6+GAz1WzBUMz91rCm2YaayU
P+hLqTJD+LuqAhs8jMteOMi4Txq+De8yqxXoIIhG4cd3Cpk1q1C0Yfy6hLdSMimQ
IoAM6Z6ZoQJOS1dLF5nDs29BBVP2Raw6KBgRrJT83qOyc3wb/uTX9fyLlAKiU9nI
/0+FESRQH/6mw51nTXLwOFDbbIX9RTHLgGCCv5HL3Gjhbjjw7zLggnBoeksgTJYs
0KET6yhI3pvr6rxelxJ44ukAk0+Mz/ckhwN5TQvsUe9oSjZJIgNmXwGW4hlsjDDI
8tmXk2ioBMoTMK68MZKzfDQUeSCzzzvAVANjr5w6JaqfCjlDgZSkGM7pL1J7G8vf
quDD6onwDnS173lSzzWwu01kTmlOWmmDIYbSfLWZexxs9LPO6VUHq+nWPXkgymGo
iJ0sYVBkjzLS45vmrBmbiirDUqbv/O3UbPt0MfLFvgI+3PsDrFKcW7vN/O2AqwJ8
UXmDj92+y0ztE0UHFddNtW51DUMuhzPCBNc34R8wEZE4q+6nVARbuzNWjfajEDd/
O0dyrVUlnmBeHTxv4RI9VdYPto2Fy9JISQEhsGSHEXRIGj7JfSpsfoAUP5J4QHWQ
VjiMvkZPGkxa3c8d26IrBQE+ifEOHjHXUBhNvXGuhVD//FgFHfKRSIzw98vinSjW
rqY3J218FOf4womojqP5JtesypxGb6Rp2uZ+CkSVrJgaQDLqP5ZwJb6uzKYuyVtZ
HuBfYjeGDOocVSMBzpxkf0sB/KsXclQEX1caaG09lW53PB15PimnBCyTKOmZlwwo
7mLiZAGuIhqrnorDA+wP/q9FWv5gOHax8Sleh60uf5789PaXGisOR+FVDExIumw0
KzekhNa3XoRaXe1dN3TwLSDn3e6oCvuRax61aD7fhttqnIYlOygEEV1vxcJ8k7xw
PLgL+RwNizyPeJJGRKZqX6x7dtX2pJwMdHoYT3xhQE6DjZ6sXx7+E1n6fPdn5wSN
fPxYauMcZePlnW0mjdTo72nyoiEcaW/+Yfi/BQbWd9aT9qcb6eS34/PDU6SGcTbi
OOCfXW6b7M2sDSrXcGRS2/rws0Zm9TnSvZp/ym5XLPzztK0vlUYUBDPFfOHVJrSM
eAcA9AZddn2l+0QNTz/+Ci66xj+I5wjjmboo2/2KuKcAcxe+uCc3AC5bz7V/+lJ6
twgUPp1AZUpH0X+m3lqd4K9lQvtntIJek1dL5tZU1pdNdFCDna2aD49/YqSIrkY1
2mYYvxL1EaPXsue3PdXRcOhLTBn8YijzqIDlRbDDLI2WFk5yweBhq4aQ3ZAgHNml
aZOuQAMXo6/ommZPVoRNaPL7YuMBJ+vBR8NBapH1ICrVMz+Nj1PWHAov4jFo2wdW
2wrRgIjmE5kae4XUKTDly8dP83evtxplfU798oFP2HGxF4xZB6zMe+4ctED+TBJO
GN3EOud8ROHpdjVFYhAhpWqU2KKSeQTnJn8zchhIQfurJr3GcAZoREx+DJm3x/A5
Oa35ShjDbfFQJ2NOcJa4ixJQxNPHcdQM6OnS0TRPXrI3vcYIx1DpY9r9mAK9uRAC
rn66JIC2NJMR90Eqvb0ub9NZoxeRnyGDY8NSFw+mMqaSXRvJ8+2f8donGnLliBWS
F0b5+4kWVZmWpd9ZQNFKS2FQL5sqDMKwCy2LoOXmJz4/wQHxdsSw0KMMeLXiXjO1
FkOUuMAJrQsixNepwssJKOIX60sWc+ZbN8ESi53ln2sqZrWa0eXivLkAX57I2p/T
UCRWg6s97IceNEypKeFCIGh5rNibQqRT7UxpIsl4x3nuyLNN662Tz63O32O0p730
Kz4oJD2KMYy7AcwxD6k4IsbcRw5F30kjAupCr0BGEJZDEGSI2qCI1W9bHDQgYrvx
7arIQq8++12Oaa20HYC8I2NnNQdRK0GqI1w/C9+077hT1+vVkQBxFuwARjywMuSt
2oBT3s9Ey5/yAZ+hFpXjlgAjzRTBzkXXj04poBl7T4JK6K5ERea8yYelZp2PceuX
DgQPQFc5Ba1fvHNPu419grgeSnB8EMpYGePei8zsKT8ux8k70v8xzixxjycb11MK
r9fo4slWjti1kKKRT1c/ACBawyhM67av+kPVecUhJhyE7sctAg/BVRPCazL4MrVe
0mDB9eLjNqrgsNk/b3/+6tUaSXRI7fKvUBdX82pAQr0+EvtxjA4SiQ0+U6NAImRw
enUpmqem4elDnYEujERDHq2RMOHGAyn63mMVf3EDCPQ3KMfxQtfP7hyuPJAee/2K
HrVubBLyB3OzGHIGJuFXzxDtszWh1nGhNyUNYNmfqzBzJgvSTva6KkG3HJzh8YLz
7kVTj8xzXmqg2JRUn61prsUqW8D2AI7eklbXcr6wA3FrkgP46QaRk9CzcIyudeQi
SputSgC4Gc/2Z1LKrsdDrpMZAeK67D9vgT1dU80XzoHuiEVcYxPEHC6BjvLNy2He
lp0c5nASRhoIpqZzWtlCXJ9B1y6+E8efgjwq7QIiv4rJb6Mkc8gtheaBTpO/U1a9
Xxy9ni9FBQW4i9COkHIwbB3UlZ4jnGdy1hObbeOMh3rG+kk4fsVmzS7S0Dar2+N9
xr6/Vm1e+tWZz/uptnk0EyP5RRg+8cAv3fgJdBHSdTfjD9thVzU3+rlurhA4lISJ
nvhzbHefoV5FPBIKxDQUXVDN1AxhtVniHXjQVdHzb+RucMibUFk5K58uxy8sMs8t
+/fKtZrYhMBq8oiJ9nVR5coivodqtz/TE3yoHfyUoTMfg3+UXfiHj4y1/QRlbDEf
nYEQMow79b9g2/Q+VeNLgP0ORPw+PCawk3v/7ODO7kX4gtip7dOXIab1qLiGAi00
Duu/q/RoLzG20+2UZVNPKTBQ41JG60vn4akM6OKaOb8D6c8ODkcyEMk6zchJWGjl
Dn2lmxvuWTR0R+hPK7dlZcc/3f3qk82g8Rd5sgX3+Re7nfmJ4bx5O9xjSwOCgv7/
qeEXPXDAtCw3OMjYKd+N+LgSGFLZCkhjuEJeNjdyhHp+3mkRsBejNklEbiWoBEzi
qmyzZbOBIKWKxO3JJ/PeYqdn86qMhqq715UdGG+z8zT3gFJVE8rvxj+rANAOJzVe
uoSgLwxocq7swe5V1KKHBzqk3734gkEk+R0ZNs04q8dtc6/QeI91FRgxUkdDosun
8ZPYxFySehckUbIRVxv2MyFf8eOp86Zw5ECdPEQCx4tyU1nVnWRUNTXNJRRc9ArC
gUbVCqf5NxF9zkfUi+AZTgPUrSYSUvOeUU4LbE6hS0nnyPunZlgMXD3HgxiNyYaA
9B2MriYpgX5pj85I+hzgztuF/hImupsAq8P08rwBe6TUyRaryDqbPp6GN+I4OneB
qCNZODMpH0QBmK1bUJk41y8KVMMonA2lSDYHbJn6iKXEMAvFPzqNi7YyA+mQA+mf
Qta+Xw9yKaopvf1HM5oYidUhdIU9rlfpzFKjiiWJQOWOkzpa4xFB8K3Z3/9Y6K69
KrkmbXseAtROiusxZ+/zgAd2VuTZIQouVrmpa4/er8T7SCOMRlqnZzoWwQ1afVzo
zbmAQPK8twpYYXmBr7ngubS4daPys/wO7qkioyX9aH0YenAXnVxYo8hz4SQpQuT7
6X20hhnrKi9RJOBiejfcBpV/RsmetshA3ZqsA3HyH/YV+SG+QJZyXsRNV6z9QYhB
hSADRYpCh5qya9QX6AQHyJl6F6lRKXLa9C37DWYy6DTucpGpWC9fvMjznIE/j/NG
fnnN+CCW0zCCgOhiblMSeVBW3JjsC/VP9PAVFyzSt/QnB6I46uufEPL6W82iWydS
hs3dkTyAX5gUyqNdUsbqg5ryeNvZiw6StB9RYBGkFxyAuEhsJJUDX4tixuN2KrZu
5AFmtyVfegOVCpRhsCF+AagH4Cilf2U9VZoN0EvPZMuxnSGuM3X/lV/wRzoKCYzp
PYtCxMsugW8UUQshRZ0cLabZzbFPwvaZYTqD0PQbsmcSGcGGgIz2sJoqLLNCILlK
GgwzpjISobxqxOawqKFiAOY+w/fwiVj7MCVXbyqYe0f304h+Lx70xIKtam3DdcgA
vnGc2D9vXUROItFHdhH28Qcy3GIoL0bOtUkZDrmw0WUjqPHnqLCbdqBHZ29gyeQP
/NUth7G5Bg9dtwnFS7KjKDpHtasMWjm/K1bLaxQzQ2xzjRZ2ddrXE9ZPYTQAIoIQ
iVOWefCiSLm32hXn47RhIYcRmkVt0U/aemvA6NFfGv+Cq5GdMYiEJF0RURndRcNg
DvU4IU0moSgDAjcS6n8f0fo+Itx0P3GFMnXv7QPlgt9k2dW4qBTIt1yW//ckVoAv
NLxPhPxlqDPpalBEZyvZEm1D7v4+nPT55WOeZXssogJCIINM2Pdvsy5hZwIOfwXK
XkY88ccNrBmCNOS/q5cf2yEabv6N4gfBcOaTlacVDtBItEWTOxuKrSHQY4HCa0jj
pRej+rcRFR94GwhfEOgAlSqOiLd7+lX9U8I8Jw/3D62PDFgn0K61Mnp2eAv0fQ27
07mcqIw/i5lxw99CdE9gOiRN06u/1q8R99NvwdIjfkP/mZ5msnA58cfSQJ2Y/nTN
C6Z2fbD95yL1jRSj+N/GPt5AS3DsQQH2J0PDt5jUkexd9pe86OAFtphutmGvbQ4d
QXm1HYK6q/e44vKF8A6BQYae0MJGW4jhmjSHR9SGLTXsyLE31mLFx+7Kc01hMZf4
bnbpDWs/kRkZFSDvr+GlqN8w/OmUD01b+xdhcortistuWxMDC2MRly866EENxPqI
MuXy1NhdHdALRUiB5qrJqmbe73T/JMPmSYnYtEtqDSauulPmyshboToT8IgQAh9R
UiJY2MlQRAG2GIhK1XQLTbl//W1zNEwOeOTmyGKNWRxQsw6Ukpo2bNiO9wGPHjVH
CJ5BoajHYRH+zaPfWyfvk29JXFQMhs8PjUwLhautQpX55rFWpH8HXxJ+ILJOSQOM
xMnEWJ/GJANJvhI6evs4w7H3lh9rxx44m6K2dGnvI7Rb0laFaTnAQwEmgYrxpwvT
SWn5tbfO7NYhY4CmGineEzvCei4+p6UJyj5P8duYYlIsUvfZz9epcybFI+Y/bw9p
RcPnW7IjMbXo3I0vRI02dIKQmKcTwTwtv4RLJg31r/s9yMc08IoRp4LenLVulzDT
Wo7TYMmuSqCO/KrMr2qgWiB7euTnLhXJepvpNedKCBoZqwWBkTwyBcnfbf6yksbe
rPE1/gC5YO5HREhxD41QBSuwMAZBkE3XUv9xP48mSfFC/EP9wWG5bh0pls3MnWNP
9suUoP6feoPg+qmKUk+YJqm4RJ6nh3CiHllIevgL8HZEBGdlTk19ccuz1J2kntpo
KC18zBGpKHwVIy2zyv8xsnWn4SJjBEhXtwQv6vj9vUa1JDpeIVsuDGkP935uqWJ7
g0sfW1xmnFp+awadRqjLax5nUDsuZ5KmemrDpbItKV4adEgiwTG9FmjMqla7q7/8
fpyfpK4IRs45a0Ur/PwQ1r+CI7RrEyNswLmCN6YahvCcHXQR4S05gUg0Ble4GjBQ
3XjzYwHOuRTOhG0SNQ7A8JdcooGpEzHDOS+pfcjf9Oy9+1yH1rJM7dMeGcrWIz9d
D5ialBTrsA9ScDQH0YPYZ3MMWqYBE4K5cWEjBpYaMR4RLBqURBLB9simFFXIFwCn
f2SJzT4iz0DlSO29mtNQMM1YSPXs+XT8OnbWG3GWTUHRoRHTWvuX2nPJiHg8Apak
5KkEQN72HqDyrDwxR7z5U9WlX/IkoRojlnqWsUyAiJ+QxBYb1SeWJniO4N3hKAbX
bjl5ytzpANoLXkdqYjOMcFZ/daTTgV6ANMg99D0tFkQeLfD+44Zx208RPevQ8AHF
2PJI6BXNOg7fREOoiF8v96xHq0itM4Qp9caefuo5KWf8RMfYa7/6xza5obYwmJ2V
2WeJYIi+vShF/Rq4+jvXUXeIpiiNzZm9GefyQAdZnnmia0SSyZvsOo7LXrEn5xau
JmBS221k0jIXL6Hf+NQFkFHLbwPtEbo4++RxZfhCwNWuT0ENThslhLbk8cfhK18e
/BQtn6/1mvrc2v4ubz4Jkk1EWvjuL4O93H3q9yOaO1Iw7RLgjM+iy/Lc4HKuDRys
Q+5yB/fYeZ/PtqnAhhpf0Iy6+VIYRc84KUJy70Ki0l605mSpx8WIhh1MVQLp5Lhz
weM16knJKOYuan0Kdl7zKILvwUdNRV7gdJrmzCRy5jS4WtKNoD/DZSjW5WLDQFN3
ksOL4DC60NLjv1aARDjIVYfke9VRJyqPdKqUohk4WU0W/dxn9hWJhGCK8+kexZWu
m5uauoflOtTyDBw1buQQcwAh0Gs1x3X/nbGAvhN7EYrBG/S83Q6hIZ61lrJBAnwl
d3r2tc1DUP+MrtVlD1Oj1popj4fDyJK6iEwNNcc5EDsXWOx5i/4EDuBSflAnD63w
nacH1iu26D5P907//NNqKbpRKFwuuoToHI9MblK3LrE3t40egUTLY9OsobGDNTcW
3EdHR2Brf0sIBxxi2O4DPsXBO4iVacaJmVOz4xQEaQeDCXe8WqSe0hivKaYl7ee7
rRlit5CLw+Xz0G+1oi9y/FjDsquMbMI5dtlSs6eGL0bfmSO0G6oTKzP7EdXg7niB
z0UYk1Q+ePGdaDKIB5Hn4D8AOIbgSel4mMTQHftDaPC1LKRWHyrGS/9py+rPML9t
rZBTDUgKHk48nKjJQfQ4rF6+UD7lH/mDJJrJbuohx+Jj9ddaZqV/Z1+6u5B5dkEi
SrnV2fO+uuwB+gYwa0/LDtDLxnsMrurE6vXEcV++pWgrJHmWRHfpGvvDpfS2aWvh
68pO1173ts8pVLgRs3nbcyoilfsO3y5FmxPKemldxZq2Em8AhMRVPf5VaXeH9UO9
9pHzToGtpduKRHprVBoiZhD+ZLLUsR47LbskTy2TIRE9UiK/S2gdKxjiNRpROwo6
uZfCwCnzyXL7w2kIUD3aYuVjw7jIMNnk7xyWgrTcaWbsUqiFBdXgqkQyT4UTBCmB
HS1TV6ugddOQJcs3mRr997IWPfAhBVeM2tfVhaI6SFS7FuBJNKjadUiu0+gMNHUO
kag6dFOQXI8QP9jtGuDIqwJvTU2lGo2jpoBWxwtlSW6vYi6ebkekaH7IAiUURTtL
vgNssUcFasPDZN3D5kFjuVUvWQqtBtRdebb5qe68EMh3Lst6KE49sdCP/yKUKlfU
aRx3/xJ639gfLbpYiNoh9qXl/Hgpcwxi7XXUGLAYtLyAUL4BaeGJWKQkXnGpDFhv
t+TXwngBqMJmj9HVK1j3LnuZfj/3NOzG7wPj3xeqYFmjAhd8RbRvRg5ipgxo4aPU
q7vkBWxyFxf66WRsYr1Hqg7LeoLzHm3Ol3AnTUtoLZ2f9jcFPLh/oQbfvsUpiRqD
tdYbYMtvj6C7W5fk3GPLnJI3FmIdajJfuTW1ZwIgTUS9zEXMhAmFNVbWv9SfAYu8
C1FovCBiGyirt5EubTQZJU00Sxlk5ckH/r9npcq9YEBXa+r6PhLyt3O7eH5mDtjR
RbjEDoCYbLKjuDOuxWC2tDzUshfHzxHfBKdz1DeYm1wKtxKkAxIQRdxBbAM6t6Jl
PDBorNXw3HotWASUIG9dq+TNIOgyG/DWV79waHca5stN437IVsVVLmiXb7lIgbus
kmdwBj7qm2Me0IYtXFzTsV+xr1/wMjx9w4+qE8mP1uXuNDoD9uAjoaYAQWXrBoWY
3015fPFZjUI/CYzWasNJ3OxuBDqwUbhmdBJc64ee2PbhYF++WqaZIgSH8+c7PURi
UtUdSAZ6RfleArqr4QlN8bJoZr98Jq951h6lWuePRzgFhFWITWPfQFAse0hiTuF9
Rl1t/3EOuNDz4lvhm0RhmArc1UiOh2bsGEGbA2lchbDy6KDn+IjPN0fZQRC7nkLk
dGtQ6Gg3dkE7svRqBTX5nYjw3ou5Waux4KdFWENPGNCGBoXuXSrAZiCi7SlOD2Bq
DPYaLwHLColI/3nOmHWuQj6MotYK9TdaRqFuCtHBBPY/rFOCqlkqYJTUb3BH/Ic2
2oTvVmjcBBB8RoKM5VKnpmYGVe1BcCpgcSax1Ol5YI+4RJCBJXuPISQb9XUq7Ebk
q5TeW/gOyQZOAs54OQeLueX8VEAx7f2h3+i/WSZ+D5howdeok37OPTisPGAmHra3
K61K7rMoAaOEU8bjsS4imj2F2Gl1fYrTgszKmyhmOQqbBxbKHq2I6IEi8Ib0QmVb
HOBl7xNBfO1CZdwRAsrIsV2OaqKNy+IXi8xht3FwfAiBiMPejUN/zT1ioCjaQTmM
RqEvjJDYFfoZ29C2UZluSBMNZiWlYFYNYbJndu2BcF7Vvw5wjWiuLW0Nl6nipZLb
n9SX4VUTOsfVKeczzPZC1BvgYvRpejvE3h8BzZMQ6sIapc868sgxwU6VbZCWvbQ6
yF0oUnG8a+CjiUVD55CBAlAttvbv9S9WG2UePGZ76LGTzX4rxa7quJL1xw7BjefY
fg4+ONnQN6LoZJgNeOqVlpTtBeVvlNU44bLryeStsZS7GnB+nifCfZGwrt9USbp5
65VSvVamXknwCu8vURTezs9jOfY4NrMdPEuSTrSjYRNlz2akgBoJC/bgW6Ff0rQZ
gGI96GwtbyiuWRp1qCsJapwC9kRC5aZHqZVCpIQOQ24dtO8QgbtnNaSdcoH3DcZf
xwbU9M2yxicYqd0Q9xWSXPgTTE4TqwrSOpHlTEr4jSMGBLrq3SmEAH3hqzqiCN1n
z4HAjCvmzESBAyvGBRXANKdglB6ZzqmTXQ4Bax/xMgJWIdK1Gli7reV9E3VA3ykM
Gi+W1MLYszYHjv61ppM96qLj0jyyi3oO+eosobV1FDt2lyPnOKbs9i0ryKnjdjfF
iSvH67KoZK64yYZjx6aQ+JwpC6Z94XApEf39z9LlS60Mfnsf6PSHwNL47poiRvN+
4DLdxd/P45LaQA6OyafHk80ZrsvFi1R5ibLoSNi0Z2m9h8+bufqfbGdQF8dNBsm0
Z6so+XbkmvVi3EgncOFFwJllphNPySFxeifuJ6QbSu9DNIKk6K8OMbXZfRWvMRSk
re5zgGVmLE0bGqSTzY6T0pIL0ej47t3kcSUvNYHramVUT3jRwtDSt656AMyMmoCE
uXtyd17L4C3SDo0rNMQHOzV6tUAIHBblfqCS4C3eBa10Yko6jBzJ8i20JugfB1SB
y/D4DoH/mIpqHMXb7k5ju7giRvjjT8vyE5A3Ue4/98dStPg6HfT6B2tNtedmoYB/
75sK2L1bBmAxJMY+qW51UBsWErRueWWx+KT3/JCqR02fErY97U0CDjgUcHm5WwqN
jTAOV6CJsj3/YG4WFYTCg2L5tc4RZHc1aLscf2zhMVbPzqx6HprGN4ZqJWs/aPBP
kzR3p2ZS4Wo5dIBXtg0OFByvxXCrVylT0Pt26pYdugLHxeIzk7AlqqbSNW4pCV2d
Pn0HIYZpgLAfGCB5b5Ou6vYi1xkvS/UKqshcJg6vcAqBRfi3Noq4DrVDMq3/AMul
lUokq4Octsy78DhfX/f0WcQMCJQvn4s6F/+RhkCEeLy7NlLHbIERfRZH77Yu50Xe
bDKo62/vXLV7Yg4NncJCnR2tKpmYVwOaD18ZuaJy+zLgUkv9CHifz6jscNfO2W/O
CvHF6OCj0Rzq0xIWZfujCxEtT3CQVL63z4TOKiQLu0TB14vLQvQfQ7YwaN7qeEQ3
EcerSzW0XZu/VWuReNiPQSb1+B5nA0K5qFSP10/kO+CLU0d1DuEac9IvAi78EOf0
R1u8hanAvvzTYWPDKB54616SBSsC87dKzU4maJ0xtMlQLf961SoRSpE1X/68m7xd
MUoMZk/NYRvXlOcKr44aid+rs4CgOpeBCa9mjkutsYihLzgGnZIDXKvDELYMmext
FvgSfMSdXItOb8EGwNlzcqT1J6ZYc3HgJzBqDcSHbThUmBo+YO8Z9i8/so58aOV5
Jb2s3B4T4ua2Arh/sQzwzkvtgvzNsVOF0wQOXIwfkqjgKTA4my9GnhWjMMeA16sT
09XuHxQk/IYs/fBxBiyIeUiyirM96Hrz94HphsX6V9GtFLIj316UMMb9Is68BQDi
VSFEI1VKvmKDvFLZMxvV0Tsst62BvzcXOlSkjH5bIAzhEq1674xqLXeiHE3HCkn0
fCP3kb9QdeoNl59p4dGcAfJrC/gVURVlFd8aKCcKGbbtvZV8RxOuYA+GdjenG6kp
NZpwV/0ndMb46ZUvxyH3aZ19pEGVIGISmbw5WSJ31ogoAkISQvfnpTS/qWq4pL/l
/WQkmxpMGpdhgeKqypQPtYn5kSxttfke8OfrAVfCHzeGes9qeIiJXl83iZCS+Voh
3NxOvdAr0j2VjUBuwblByaYtRKQ18CQmWE/GbwH3kdpPCbMrbHfa2eRvVlIv0hIt
0FO+NO8NbDF1ziBgp5ghN1QUKUPD87CpKriT4USH9S69GvXRHFlQsPerxhIK/9rH
lMfHZwlNepfwZLVfzNaH8zyZXSpAYQSTYMUoD3rzIrcLVYjpCY5ga9jh+vZqz7Dn
bNSDKiqdknVgRHuz0TrYgW4SjnChylP+/JvAvEnEj7hIbB5f/HEgBZ8X1mk8Sbu/
6CITAB/z4rHA1AohTdt7FLVUiJJtqYX4GVzJdDYNGWLx7KE2x+IOCJe8TdwDW1SV
LRwMbRN1Um/okv6mxLwW/KwRaUYXw6Ef8usv4VGm2UNuE5AIwnvmEjPdUF1VZo4N
AsCaycZlCWIDxxx5+WMs1MzqfXxMCtLwbZ1eJ35JsbaTbH3zx3JPZHnW7EdbO705
CuIAQbLYDSsU/jcMOU1geAXlzmbiCn5RYNS3GZcXZeRh2e3w+k9l0nf1x8eSA8bT
cQYvlWgxJBd0ZQb0niDZI/7Z+eZHBRszIeZOGCdbfoKbXLSPaNzuJSn8ZcBHGL02
2F6o2+1ZJgfBYJllsJ7oxO5Bv+5rnjYu280EqAmd3N5jbxxvksfjxojkcrgcqkbR
scmJxdef35zoGzDDFE/wdrmRtm+7TEZs34Y1+lHCwEWmLgEvtUT0+6YlRRr/8IVo
A07gUlaf3JtLj9faxEgEJTEPpCuuotTdkFyUXff+z5Ubf9D6ODcZAZmL4sJWqSRr
BsWw5pIHdnY1TCfTbZRNWKd0NB6XU0i5wq0MMadVw9AjhOySjljbFMfuR8k0V7we
x3plRqPHgi5jKDD065vyY/H2xxcMmCwim779eFvw0O7FurOW0ARHAxL5Sm1yHMrf
PcVKc563FGwxSZ55jbm7XvhrrTiYqVuj7y+KMrQLd2SryW0mRWq7f/F2ywMpEbhO
rlD7iBbyEe3Dlg2Bj8xwNyoiyl16ka4kaHbqFfzMSBOS516Z65SgGmTMjgCd9nPe
gl87OUg30sxDwBRxkOltSq4PGQc0BX3FCrCvpVCPrf+zG6pkeBqw+q8UXWA1JBWV
P037E0xITlQeGPsULysEX552OGigardaK4lBA7OpGoduQmtOylWCGHKGhnxRiWgz
Og6vvZCiu6ADOrAlV88ETLR8sppABCx/cLq/E6v74U4VLN9da+7fwfz2KZ6uNAep
zFsV8PvBNpEkWdiOl1R2HbKtkxY7gfLT4yjfTWHJL1gjjpYRK63dyGUV88BBW2vb
b3cxZp2okNbWdA5zgXldMymgTVEblN3B5uDnOwNxOsyGNGQ6M/SMjh2kHvXvwRcQ
Ancq6MfWVzpfzM6wJ8/eRq+XDqSq356ALkr5hPSMC1v/GwLr6ZuyPG7s1hISbugx
EmlThl9siYZ7mwNXgHseHYROs3sIjTtXHCoB1gmEwWmFYoH/Jqka//V8+4xbvfbZ
IXkjNoh8UuNylhfDP/o5+6QGIGXrmfsuHQcXcAcebLf8hsv7YK8v2KVesB/ryUp9
rDOOfTRchWa6/zT0dCGrcNhz6OZc1akzwoOVzLhye9FpN+FEqK6P0QICNw8pDy4S
oiV1wCSvO3AsgflzwRY1JaD9rFHrGEwUIKkJGbS+fJ1CSdtj7sHwoduUrvTLoptb
yK/qNBP/0iXNUKtulCag3iacy0xVkLVu4dLi7UcqzlSYXtBKdP5Fb9fznU4fvyIA
RUBHeDeeBuWJrnBoGBOnP4HKMSsAxamt1W7Tkcu2uzb074XeCL22elhkKF8vF0jr
OT4W1DPV885y0+lehY+OGS9Y5sp6Q1AjHfEd2OqArtbgC0lw0LKcVLYfb7x6cA17
BK9WxJ7YMWL1/OUSWVBdSRpfLEFoeIIiY0SZvGXIJ+l0J5ejBXcvsu9HkVPqNGl0
5jZV2ATp94GepFRBaNLG0Z6IeR/7+SAMX7AXAFRxvdaRybcWnF47EiWP3Qvtce/J
6p2QPjEBEoTjXbsO7xIaDoHnAzQX2gwUAgw3mrxFqGjWrxdRr/2RsEGXykSnrFCC
Kf3oZh5dtbx+iSxwy4GP25N/b0Sw2Ki7kDfJc5BWSd66UKFC8YDg/mZvvnfWwS16
8YtFa2TK7BbKdTegTFx4AXyOj6HIfiarfpt7sU2jTl/++MlXExtzZlXf+WCY6bbi
+HB79rHsgv0bk+pYf7pnbC1K/VS4UkbQlCoJUDQFNDHklPagP/I488n/E2EIyU/f
OlJSRtJuNF4yUA0tx41jKgKXDp9R/RM15DhswnorG1MT8YpzXA7PxM+IvXuZA4zb
6DSIxDs4ZWAYkqNsn8ASiCdvjvXsVJhcENLXMCmwKqQTXR8K2Wo0Z92PSiWC2nBa
A4zyOgggbzUTowCjDasOmvOuucZx1py09KP7c3wn/jqUZwbmIrTaXzmTE3INNPnt
kubd27POfbtrLFw2DcYSJhVpWg/bvz9+Sid7PKwcLolBcEd5CYyMgrwLBclZ60MN
YjUlFSD1W+jVEsmq9dh7cNZD8uXOU+TDTie7pNuuJqxrT4Kuhfe6uTI9GckJehaH
PZ8bOAG4QMozvU67tDkRgfzNxxMeX5xtRxHBGnJAqOlkK4nyhr2zOATq/Tb6O1cs
NmLeuKqU4mbNQMVhjRTq13BFk6ZN3jSlL+5qbgJzNCE3ufTlW5co/NXEa86r1pjm
RoKlr3odmapy2/+89B5HWVLicMGfp3qi26ENJT1wo2iI1STDvBQ86Wpawa1txw4f
YDC4eownpYsrSCNvHavLplcFFiETqwXjOT+rXyBcK3mYTfZun8MUvxHbEpG9As6b
tN/NH8LZjFHjPi+QHVfb4cKQVoZGAoCj5z/cghZviebJWUpAHcdjMFRM5ZdGxD7s
uSEvFWzzUNpy5eZLrqFOMpaNvwFct6Q0qnA0tnmhSsaswDmUs8Z4CZz2W2zINLVz
eWlarLcSHbxoH4dLtF8EaZuO+krY86vqc8OemdvZ1m13t4dzclvqjbBqLp53kv5v
uU7KMTtdytXqId78My9sVGuM0cXf00lIU9uZhZwcBzAM4M5lpIFxx3zpQ/92z7F5
S2YI3j73MDItpXI8JI3dt1K7gMr89+sXFUKIKiEIgIynXlux5vjFjvSUe0Poxvec
zDfofxzp3WdkfjIh8gWJtv+QvGf4wTiAycxku2JWOeknJe+G9Xj/N/ak6Q2ed8cp
xMwailRE7VoBCcjrZHctCnLak6Enl61JIV2UD/59ANJc/G9tEVHMXIFbPaegypfH
tnvOyQ7r0OQT3Cf+i4oCzCpfUluBZnClA0xu2kJMirBcJkZ9ImHgk2Kcr3W7B2a8
D0Jg69iJrm9esmGuCl3Wasz4Ee1jO/7Qrh9PNDBECqJTDLCXM7hlxVlsn5d2s5mK
k2MzKZa8hnzcvA1F95s/0x3q4TWRZsg6qrqaQO1Iy3ZRbj+zYvHMjikS+3y8/MhL
bjUCjl/h51XIMdXVUuj45HyBeKVY24HKlMLl7H7+w3t9tQ1AWkMBfGJVTb3QQfJq
cmrF+t4tNuxnm8g7xM9ifM4eJ0OFaqdbrLiKxkwXaKm43quQAEpDTndhPMCHSw+p
G7/n9LoyJ6r5Dala4qX6YCcXxcOCAGcej9E9pni5W/onMTOJPBkvol5o+D4DdB7G
p0vVoCsVDfj/oimnuXmLmTliByArx1RTu1tQZVpNProQBFDoFB/71U3TGPrz1B5p
mdK+vsvOlVajKhlLZZuB93vX6w5kOX3uboNQzV6vIXwMjWkP1aFiIk3Si9xblzKf
AJLPmHBgHa1XfcBkqzXjmqbdY4LQvqtSZNNGfufRLdS/+0iIEy99Y8xWh24kL1p/
DJEtZiLrX/i7g0cD8w3UKu3yP+NHa/8mTcOBeGt1Zv7pOsiMvAHNAEUvKM0dRB7e
Zo2Xf7FWsVSxEF6pYH9o48q56r5qAYnfh7lAh9akNcAPJep1RQRYL38bT3BS1Y1t
Y59SeBCJ/mjCLvk+yIUA1DHdYceT967hPx7MUek3vyy181iiKw6ddHeLoL3vnFJf
iXIWERJo0Au8wd9kio9JzwyG1aJ+FvaWXDUwJxqHqJtmobMYfXUVmdrjo2RUPIu4
5gnLp6pdnv/zVgG3ZPnUFQ9qv4C9bXZbSBFR9GJOFGhwEPzu9S4FJ/7stG2a6/Pl
CH1kqjYPHS3ehsLXd6Q8rpQVkpBGdYb608K5TLDqVl1Pk42kemVrlNPa6h+YGeEY
aVJtIdMXl/yH4oJDsBYu1NN7iThRuBpB0/8Arpcr6ODrlLfG010RYB5rC7tUQOEz
4ewtT7sOFuYYaMN904TRJG/H/cyqyfBRIJPK+naVSnI4omnMszExu0iE7nxZmwpT
eONeao7FLnmXoTJqJVBypWxTijp+h2dHhKX6XMXnz0oHuK0QgX3hnzTKqsZIOCjl
EJZHsVl2hgyRELDdHLGe64YoLwEsz/BZDflAY5ynk5DIgBx4cJjVpYnYH79560fd
RALJK6bDFv3rQKhXWTeLV3gD+PjtxWZ9x3OCWFiVyW5GcffNz8CLpjS/W31Iolon
6pWGVeTocFyfVcUB91gylYdz8qUNmmczjxt+6GINWDn1uI5XVPrjlplAYiFC//ML
G1pBw2Z9Ppo+Xhi2sIBvDGGNsrh3zeHQoVv0Cl+rfR+JHLyLFvMAh32xpA2xZeRO
8DLoJWvLfgkUIKxN2e8AO9ALlYH2z1m3KCEgG+srNUEqlqsINtdoSYEvuIUSsbW6
rGHY3eU+yHZhR+6tzJ37rF11qQllvXQB1vIhPG9UhCSoACJByg77Z+I7qRRqZrza
B+fsXAPI9umL05+fy1MjBXTLibIKHdlmOzwmNFNma5k0sCo1oiHhVnaor+JYJqjF
86cUtykTkf++VkD6fTpOhcQPgdMHMYvuys/dlGbsemHJSwN21EFFzpPOsWtfu987
BqOTlqgpKxTDPSjLNXsqnI9ry7L4pGWsDE9xFeXYOzAloU2S4/K6Eu8JAOq5AZci
34H1rc+PabyaRR1Np+Dn1L6vZp0ZT1Fp0jCoqrNi1Lq+AFzSjdofsYWLTy7iVVCC
gozT24HvlLOsMz4uheFgGWOWp8mvVIQELjUJ7NGnVugwYarCFF2Rj59jHPGETZvK
bRv8wsJoKhin/KeWm8/DsaKZXOYWm+bRFJ71gARxkY56wqrUZxzj9YirUMCEiasp
HHhQ9EfLGWFU3XNZvPB7ch0culaaDxy7pmCZw270G4YZw3LMylcq64GIY3+MO2Ss
ldyhFyIsUmoxTY/uFdKSkU/xpIWvoeIx5Gz37tSPXMVa5OGkmLkr2NgbnL8G+wf+
dGa1jGE9aNnWLscJ6s96YsIzOEITxynIgy4ATltUK0Z5GBT3UXX5+JeOPsq7Vo/D
ZxBsuzgtdPLcA8C9B0WvLNuis8K92x7I9YHb2+tZBIwmj00t7Fg7fw8ZEeyqYKD0
A0iT5yzAj6jRtfo3WT7JwOQAmwoKpJDwgLDIbas1YKCUdedbsQdguJQnlINycSek
i839qFdW/I2dASuDC8C+7WYrzUs/vvEWzB8hT5kvMzVEf6M/TUj5WfRUrbrfMIZc
mJeTm4jk1ZRq8CKhzcfllJLNEqzqZ74VbdaRuq5KrIaN1qQd1vnXhm97ZiwXQjJR
lFsT+nf+RzZgbM/FEWa/O4cxFD8obm8LL3LNW7dvcKfma236JIA3lgAhDhzNswxS
qseYcCN6BKHpUdNbtsTkAv+q2tc9ho4RJQImZUilZqTgo6avO7pJKAASXm3tqGDc
EdcWnViEL0BpoCJsxswNFaVl4O45xNksnDtuFwGU2ACExkPZHKdV138u/rhO1ozl
g3F/9w4fgYWhoJIyFZZC6vmvsgRRiBJhsORCOOoB/XrIFj/UFsXaYQsirleFmX8n
9bK4wg2Y8eBOhsoJpNM85fiWfouvxp15oYMiXsxkR3Ol9/GSmz6zbAel4jOL6Rbz
SkhGn5gX+bEM1LjbqPRLLSFoy+lXORseqtC89541eonpLRHxCoZyMKub07gFdmJq
zFA+C6m4VNtHnX5IJdYT3hAksEeehthPUYXponbE2KHm/NwQjokwX4YByF4B4XAf
VW4MrzQ0mNCOIYKF/B6vVydtnnSpNImV6A9rbzxyZ4yfKkJjlmWlbQ+1uX61EIQi
sCyuHpzp8obC9ch/EjI8qNuvhh4uiah1vpgqyPEtXWSeAZpyLrs+/EA4dkCGEr62
hVM0xHD+vixJmkW7lWfvzW8848B0nTyJocj52zo0Yt2Ex+WEP+skTfChytwb66XG
thW2cS6IiQ3EFyxNo/2RzMwfyUhS2vQY6hXDs0lH4u1LKhodokv+WICeO53J2mLK
ovKeuQ0S1Dy0SGL6qhiFUrz2NjLDxSJ16FOJmjvPh3Ql6tbiUf5WUs622Niw1Yny
1Syd0uep1ruAQITtDOqoQUDh8X/vec8R9TdW7B861Ue3JVl2zb1D7C1cV4MAD9AR
8FRPFtmHR0doLnpN5ZjlOFANceVU0CbO/8wOsyXahJT99qjv1IilJ2xz86rms3vt
fG2l4CueohTpmUDLCLP3Bdt6U/JdBg871tNFjoACM3mb5ExbYGrIcmK+oo7IE7Jg
G4IfzWEvUILgMubx/rQL4DV1iMP6LH7MbA/I0TFWKWy6XES1WPb2t/6mQOeQiXhg
r5uAyc3FqsFxX/XuLJYsdAi7F31F7K743BsgMzP9IPF4adC/lYTJQfbibCaREIBC
dXq3JbK+UHm5G6/GNvsy+s//FwF4nU33j+mvImx9888wKLBfYkjoU5bvH0JIWJnj
c0QdP5CHMi2koBDxQABliXDgVgWi8FH2lAadspPMmn3ggxH9XXbsyIorvPplhx3l
Zy5ry+6M//CR76w6vbwzr/qJgdIHKtYb03wsNDGoH66VCi8dehLbDI/DnAWxeyKG
Ipp8AQRnSwwcyuGGITChHMru6IMBOfJvp1QUF3HSH8w+NgnJ1lXEqYIhTzN7rGqJ
QYfyVKzXxZ7hEs6VcWOmjXWNXRaeZ/uzjGJSY4vMc6eDR4umTRoGBtCYmnhSp52U
/LzMxuwh9c3EsdU9dl8rBCudCg+1mczQha4axAoilmtvk0mkCpMVK+3eICiU9AA0
OT+eq5dWbRQrsYvcB7nNiaXVmQpMjJG8WDHZzXSo62VPt6Je2Uscpj7IfH79bwaw
YVqf8S+730vMQvhHzxzyFmeSRczEMZe3Zc3JaQQMSJKAoc5JZSb4HSKTALj6Efmk
Dmdsh9L4uLZ3HA6Sw11WBLZUR4UslpMLssIUpbmWaw5B177vMxt3QX6h/4OaIE4L
e7kbrGXm8uSI1uRKFB7Mucz8NNzqDTBMNSxhYYIHA2dUUz1/+UAI1tdvAoeoJanp
2ZFKTvT19/a0YVBOVCaJkuB4YKLXe5KhYGQzSUHw43SR6npTlw1b0Jsm4GfWvzB7
6ePmI2G0VfdMZj2sgPHL5htNdA7vw3RMTaPJF4qYJjkdD+YOU9Z9/8QFslcLFrR6
ck863qK3E6Z6KR7i66Wnh7V58os8fmddOSLFRzTmd46v+vMzWY0HGtXpxFwT4ym9
rPryvnFORDBrhMl5CGSe1bS0CirV/4bPWS1Igdg71+uZ8EUWa+AnuVB+H3foRTrP
gdQZvqluRcVTVxBE+RAA3IXobvbWF7TMgIGhJNJfvKC062QhXM1xiZnBzObdXTxA
nTT9PG5Q1w3cs9hYbAJaUonxr9webGNiB66fCLuUWh7E0QsJqh7z1ia3d1oGXxEy
g/Zl7Om0Y6/7sKyewXv4OLnamVFB3xvKUiZNxoPFcgu6z0fgAw7k/mSd4qZz/6zT
SSwF8MIpjxVDR06Mncr3MyUNVZDRDUtAfLcSq0kqAVcrQePRqSZXw280hxeLZNhn
ef0O10XeY+TUI+fh5Opdb59ndaqKTEQjXM+bnrP31uPySUmMkkGeD8RkWSAQkxox
rrpWOMU5ZhrKbVkmsM82eGvW6lqBy2Xmxb/03su6CjN1x2c61nViL+iiA2bayxF4
ZJNlZzYlOn7zlLlaJ8NBbnRVsSDtuyrqEWb36jK3+s2q73H/rY7WuOLUV+ybDWSF
hnvpML6lq1imhGeE4ozXixF/cpKHdMVB2tSBtKHhFfaw9+nLrpOCbwV3tzLrGDSl
Y2GLGnOxeVcEpilPk22Ev2aSO2Bt3PKvPsHtzKN37Oqzxg+n1Q3PKbsf0QlklGob
vHJK9ssGL2joQrrdszKHx3BH3hldIGwNvkPoli8qIn9r89sZjpzyDh/e+Qf5RdIv
Jnw4N7+MP1ykjuhnn+LcaHcS/GLzLaXcyMHq1pPrDrhZQuuM0biqVMx3YGojS+Ld
5N/jmufSJwFPT6d5TVm9lZUiN+6UyYtISoiv/ys3g+JuNHrGk/GA6CO+jfMD0MYq
S+bqlLaZMakI4SfgPaKTDL75URQVALH0qI8Urb505VWDXwwSosCLbfkSIduDx+L3
YE6Ae/BnxDRjNN6SYl8p7NFeXpA80f+gBew/LzQAgFPOvIZV8i151h1rjXUSK3zl
ApE4/zxWsMYwNBkYkmN52u/GKbTkXZZ7fgwdOcStKQWu6mxG4ZgDChIpk0LBVGyA
Rokn2vte4/SsXmk/HI3630/8NkflVwLsvNP7359flibGeXEehBX8CnBNYP3MD1rP
jqrxIiRoi3GXB9+Dw2LWPDyVV7g0eLpA0Nz5ZCBUcBPDhtlAr1O1mXcl5GMCL2SH
+nXwTEec90uksKwrUpB12/C5/kiVxCXbqnIEKmJgMkip8VvNB8KMRIQqyUxjMFeS
iHpdqxWU3M7EY69GBxQiIxMgJO2PvrfGYFpipbFN0vrUbhjHDu9y4b2LvPzGR8GR
DCM4LSSVKr/7XXcnB5JgRTMv+rXFyVkR1tyRgb+vW+2LqO7tjXtfqiWvQpA+cY9l
CQqGZevVEITj6Rr3hdeKWQWNPyjFIH49hbsXfz0mcvf6FMj0/085zaapC/qYuLQj
uqrWAbNhD1ux5TDp7Q0FprOFjvsrhExncjh9j1OhTjBW/p1pVKk2VGbpe4GfYB+0
ipsM5YEwJNunpKVINHl0grNpqNYsJ6BPqG/Yz3AhGLIIfX/LbNmgEzZUwgttP9Fx
Sk0UF0XK8Pewxyz8wbwXDyvJ8gCtPDPeTtrmHPieonCX/g8xWY+upyHSacG7fjh6
ndzs57gG6ql62ohLhTSwXDl5uLRSK7SfcwCjJy6TGgF2W1RERULRJFPZp8b/3Gyd
rZcqJVVJC1nIYTuSbaSVcPVF2P79B6iYeiOVP+Rd7luDAWcSYaeONZJhXn9/mxUj
laq/wDRdhmRbyEmUdeF8gvpdQ1Q3D/XJ+vvzodeqE8SqXbjvD0MnPcE65CplAuks
2l8BmRigK2nS4wjgNrsGH9dDumdPrbSfe3bg3F2EkJG7RKyNetsq2IEJy9Uak/To
mBne+9Lkt6MKMpeB/PxWXGxZ1JFmqdVB2K+qUb5wA5V651JYffQYDwvoccBPG5XV
VXToYlZFLCAud7wCEWXoREz05BJzJwBtGK6g0ePbYQ+WBGF+0Zn4lUlTNtij0o6s
Ho5frD5a+GnsM9lDNOF8b3T9Ffy8HK5hi/NADm7G4muN7PlCvNO5uqnCKiN0deyZ
HABeRlUziZgBxIP2MKv1esuIhvk/7t9t6PoL9zu+bXdaDSFcptcGKhORcQZWsEQY
hba1fRUcI/fnI+Q1J5W5gpeTbO4n48EAkBXfydz8Jb/4e+ODZSO1pTt9Xx3Dkr7h
NP9/uYWJ5b7NIV8uKBh8qal+o0FOyMYwxkUQiTjgeziK9qWHy5QpieavKrTCmlpx
YAfTvhBIGlqRNx0S2k8p3w3YWu70ds8V/poLUGHBu/j06o0DJyHvIBppHyUVsOPn
Y37WN/fxsFNEIED5PUNwovejrK82nxEjVo+MLoo0z3k89/cGIZNPmwMaXT3fntvp
zUsrYUzEkjeQ0DAqZlytObsXmBgy86r3dJwML/g0RKjPITztE6UIwGOOwalqZXdu
U/tGHxtTt6dRbNb1UitA25pngLamqewTnYNwoVpiR5w1ZNkUDPo8X67bQGl2MUBE
VsQLGhg4C1iTbeqobQu6kDvmRQ3jpOOh+olWJmCXjTp1xrLXSumn5I8t/4hinI88
6v95b/TG+N86sPmuDax3GwTxWlnH11HfjEogpQ8eHyjjlDXyAzpsqfBr1Dnl4LmU
c1KwWFPkbd4N/OiSctqpSpqTgV6UPfDsSpG3AXVvzneGXmPtY8Q70rJYPDgO6Tq8
c9lxvZSBUZmFgnFt+SKqrryvm63R6dE29XJwNNsk26E8b4oxkTff15q5jdKslKAa
r1WOezvRhI3QJXxREpPEpLyrb00cDiJzzdwfYLEYJ0VQ4VCEN56gf9S/Yeskz/Ws
EcQHT8T8vTGM6QKBl3Ajt+H6eKizFGvgcedTdGN4kqRO+taz9LyuJB/FMyKOCStF
vc33280KMagiub7qmkdOHVNwgROc0GHAL+wVJYy2+/TDARFbWjGnTdFxBvxvujxt
enpSod4grH9p1xI9z/CpLG2o6YNfSaG2E8P5LGRBLBKfLv7X3QPDxKEQCn3gN4hw
8BUosbvH7UKaq4x7H8pCsZaPSU+bPHJ4K+HizkTkl31dssFuq2i6P3UyCJ9JRsXj
+1opiDHJB2GCKGGH5WHIi1JlRVeoMxMgYlkZxjV0ZqMR/0wCzQqdXJIvZ6Zn7ELG
s0ILOGBaesU10W2Sl237aTrf+a64JDE+Q5VAA6W6L6xnnnc45a63FZ5eFYmjG5Jr
t0lgMTTFK9a65STSFqXPAQJFzbAc8oMIBMgDvfH2fc/WgvYxEOSM87fULLhat76i
09TaGFIIV9WJwkzZHPMAh0V5C/L+UyLx+IROHBjttAUsv+4Wcy3fTmicfyC4BGwL
sPjqtoB2xdqKi9Fc2FU7au3oQpySa1rpMQjvckd9any6mtchLPqJeoIro9wKwoPf
P0uz/kmOh2LCPw0K5YHZ1kSxHhcG7DIlDwUzCWytEMPf9dsiZEpDufwRkF4lZ7io
sdQs5zYODf9dfqMMOUqWnC/4WQNX9GwliWfwEodKr1ALdfcRml4wDRyiKLnHQlZ8
IWzTHY9438CEVK0bDyW72KjG17enRNdUxEh0iCb/fK9LqrU+qPL2zLT6V5NLdJRe
Lj3wBMb/gCoJjgSStxV6dP3f51+DZ1E7/2XSpjYQCibQuQbTcT5YocjI388jcIC8
h9kQQd0drwBuKlcUaD6wzYrSM1nPgPsLv3nctX6TB0NKDI6TY/bQNfFM0hN3D0oh
gGfOaqfPxoieNEre2rVekQUzy6pAskqRd5cam8fMziLx5jiItW/mYGTTtjAwOnww
XsXide+67GgqDIMzH49i/kjRPHkpLb6EhqtjCF/pYg+D1hBV38WWVuPXBNzQuCtZ
WycXEbrxQAiu25nSOsgGPU9UUtH27Y0FNccUjxUEhPXcmKlKVvyfmRxGsgDSKCIC
NMuGHKSwSpwYxkHn4ZFOyiTA4pqSAA2T0AybcUBhpwMwIn/h6EBxob3nB6KE83mU
YpbXbgfVMSNgKr3gahkXEn6h1w8MuM+Mq8FnYONbMvWZqEyUX+5MnFsdML4w5mYM
/xvguNpK55uhGbRYQc2hgUBDOw6cR1bO9ci8WbhU3oPdte6cjumo58t7GEKvNkuI
AmLSsa/QlvFSLpyOtZjDGCI/3a0wWqcXutpAwdBvsEUQhEdqu8CCMGbkdDXLEdwh
AzwuzIpHmvzzwm0T9G9spBzxbBnCk6ZTp+wE6NmoKv10F7rB2rIPksnqgZgkqatu
1rY5JGrMjlAM8hDtBaHhrT7siUYiEfgS+hlLfg0aNtW2eGwfKym8QkiKu46bGnm/
EHA8LXkxvAifsNU3utAQb1OHFEw38pImZGJgYH1l5Lw03G4/WmjjqgbcB6e6E12m
QeNOVv0BzvNWdYX88qB7v9AI07g+854pjFEuHLAlihSxwO0dJ8TDjDTawgYkkowO
pawOeiyXECmpExhL6v0Cn81CzBLUmy5wFCAf3fAPjhrmzBAmJWYzlRfqgS9VZbzg
BeoAXsHJ+l79yxWorO4/na++VlqJswZU3vGwAliqpYwYNPUde4rxRB0pmbuJiJuc
W/LTK5z1/UkMJ2mdnugn+AawUMrXfboGAKM0rRURiHKfQraPn3AaDWy7v3cCvwf0
M4eRDDebnnFJ7zb+UdXj4EONdiJ+ivaCO6zwRL7BhrMVACv843WzFV6sJSVLZweo
4YbUSDOddVn4Ly5PElwuedELYYE5ubBmi+hOvKbJYuAIR5iRqFn5T+stgKfSAzge
nVIrmj4uwyNSg7oRhwhpLY372v6+guB4u/EPIt8DRBqy6wiRmHPAkHfSNYHxuBIS
N5T4SSPNAaIKZe3WW2GNEdfUUWz8ZxIO1NQh2gA9eI8M9zxi+UQVrimF34DxMcoz
K94Mv4yMElUTUIOnXk0KXdTvliRiXg56TDrESjq1dfQaT3Hyw+YSwMuIjO8qEvYR
8Yi5kGzRro+0+XsGPxp7kCzGAYV88WyEa2+4I8llIG3tQ6Qp8VhyVAyq5FjnkvEG
Rh+2lT9SdYxr+MIPDUjfCfJnqkE0R5napUXSLSzR0oRwf9dMnDvMd3OaOR87eVYu
Tr7KTwDtqWqU7+zxkgs3UmWSq90V5JUfHY//QCJQOEgbak4Aj/enZyS93ynPjZcm
TIlmYjxdQLLXJlDIjjdJPIgJfIKeagKNL876GAV9eIgaS1T6/QNc5T7barEiIc71
4LifaqzOz2F9ST4j3zqz91BryBiK3cYALkTR62eMPDXsOFLUvc2ZQ5d3bY827f5z
qRMQ5q5YuLmulO64W/DTqywWsZX/afsCgzpjERgE/FwRAfWBbWmRkHrEk4qJsY4N
F1WB+EAw+dWUiLPGybxSjHOZVWpbUPDhRn1mbLxKjSh/3e8cVXafUJxVbAnzpb3I
33adfjlEl+1T1/SnM9ol6YE2M/7DmODYuIes2dWgkHAuvsxUXOVODiJNU8y8rAyD
H8ZtHccXwEmpWZEjtxeuCNz4fXgJu8xUW26j6ClfON/VYpx7TRWpX5NL5DdS5yOD
nBNrRj6gV6e0ZxzB1w4ARe+8tINe7GzSgZDNdXpqXBkvkq5hWanqNVtdQOv1bItY
SDM5RhXYRsoz089eb+oIOL+p6iw2PssxTULDD8pNyXhOgX16C34HMOxhvg0Wzhy+
FKlrN2NLynu92oiKkGtBY8lgzNqUtE1t8C1HkLcJua727lBi6taTE6NlIM8IugnF
aAnAx1ujFFf/GskWbDBNGl5cEhCyPl9dbEZJ8P2/M56VrtfjPMKiQDIzay0CUnJ9
NYtF7g479ITlbF4dmYG9QUugeiq9U4RAQYcOlIs9YwThgBMmYBsFOy3fas/feKjO
+9eBwNdNiKJV3luuk7La14kEBm6v70lMoStnb9iLpUE1tON/07gXrii5IF/nkRUf
DWAkIuyrNYsgUyo2B7JltvJHVONrm6yjkFJBXlup9hdr0Qy6bVM7SgtL9ppgaj5V
WO8VDepgq4ILdfqMyItuHCVvQ6qbAeW0p+SN8RJz37UAidKYqhGgUIHH2KDyJ3kC
esG8h4MyNsTmY7jctqkQReL/vNuie/3Obk7m77r4tsOy+Uq1pOyppwXZYssqf+58
k/sEsRic9HSjhXTungvCRzVGPnUiFYw2+WlpCxZQbrXuyfWWHT6RYcovdyrtQlGw
k1JYWd4Ph8PLZ9+ZPvXnXYvOsC+WaQpP6AcAYmj3dITMAXnGDZN95Eu0rPz+KJW5
uUxqh8b6n2jMBCg4wV4MIwnpMHhJcVds1r5Vdk+VIfxVJDclSUnXd/GEaPqQNlOT
PGs2oZCV83TCUw8rk7w8yfLcYNvYsORyGBcFwd51TEDosumiKgfXyLuNe2z4Nd5q
m7BnNeJ2uG7htRkqAGF5ossWWfBIcPrhAo1PsZQCZUCM1skJYicqMhX93+tGV/tX
dlqlrCRLQLWE417P4O0f27VxPMHSmsdmyrjFmatE2aqQuPtnjIG+d2fj37mxyz28
cYfu5uKENDs52o2z6rKA5NjsrtK6FYbaBfE67K6EZtBZteTgAs1/gHS0dI0AH/wh
OyArgQBUQVQu5wEomj4PAtnzYtRb6sSwxgKrABhwYnhHBOQjCmXdH6JiyePwONbh
mV72G9/sOTfWL6wrBaF6Td/gJrULj75VD7Ju4aZRzYjJn+VL6H7+g/FvW8Y5tcxA
UHrzOq0Q/xmojKPbQr6N8kK3mx6sOJ6h/6ngCEphO2ugHSY+Jbk0v8sPKASE66gu
NzcVQ8i/Ieig2+1DIcUMR2WAtCHVMKeI3lVseFj3nyTP3EBaZCkqm5q6VTgTMrc/
X9QCmxfbfZM7AnZEKz4JTBn6MUnDs0xP3xHT55zkQzbhFESASvjbcRMhKgxJVsyH
wNT1J6XIPTlyScrvCu9/qSZEXGVefNA0aR2F/3sQ/9Paf7OY5FfFg05bn75ObM5h
U8DVGKzXvcmIlwH3JWf7N5XJyvSqclxQa9GwG6sKbPldAwom+zMC+O0wy78jDyGJ
4v2RvP6cd8r2M1POHeCJep7TnBQuYFBKwEU4stPcezOvHVShGQjem2RIO6vqY0s4
9zKBoodiDQKvSXiBKwTX6FDXoqQMcRGr6buYT5ZEhH0lRwfPYVcvEQhAipT704B6
sMLW91WMI4MiDHvAsfhOQDhQpXT0bHqSECujBmBPw1INQBJDmZHoQIR4lHj95kH1
4LMGXSkS1GwFQez5elAZ1a+QLbxmOHgqQjRXRwRDsNWtpfQpKmaxuZd6AWyGVFNF
yw5EBzSNjRNA2z3MvgE8vMgx77jXVfm+Q8Op5BqbrW6JFpM86NEZv6TKQvLCyExo
YTjp40AeS9xcNusYiM13naApLxeu12xUbkbxSWH3bVa9k9Mbv+BSYlifytPKf6PI
xmeOkJmrwMM8Ghfsbw6JfIY8UTBTKx9cOkwNBrU9Nfi0CMqySpR5gAPPSgeL3PDl
VPSeB2+XyaGh4UzS5HaHSM+MLoJdSlSwLhzZX6mQaqcKyCBVTUIZF1OduKFAKOH5
xz8k4tZwS0gx7mNMBYxCLdxBAJyHMv78y2jyUqrxDyov/51A0YdhwmNvx92mpfCB
lsvVcMHmKLSCYzF82QK2S2SWkvPYIMDvHdYNsULk3ClM0L40+1UxQuluvcFCjf4y
eVETDzbQYjn0m+YdsV73a9KEwRoSbd+3Xfe2Dt0N3E7D+5JqwBAa6Aoq28CPR0Kd
6bEVwSH2zoN4+gE5o7uwNDxNuQXqYJ7URL7Hvi8O2WhyKiiDCvPCSjVvijjLUf8Y
ku+Rzoq+IBpcMtIl7eb5efR1xcoqRgSeOX6AybUCfDUsPHoYNklidfxIgFiVGdWQ
a3ST6Ww+NIFQcu+EkO+Ap87JMuZ2Ph72NwrTMkiRl6rnzuXFtU1uJ3nOHyjB5hBj
wrhVvcNdhkKzAghfELSNTQz17dWxil7rMUBRarPDGuUzTwJGDv86HBHigl0ePJ6o
Kgz39ndb8FlLS4Z/fbrE99gnpeDqcbfx/e3F80HUngpMIjv8YDGNG1fH37MA/tA7
oJGhQqGvS3ds0xqKzvJHV8t0tOXBc0/+YPB6wpWSlTxyf4D1Hp4QTKax/TQ3TbvE
o8VqewSRyMu3MxeBKlXE5fYVf/UuOJGK1iO0mU/H6o3wE2zsRxqg2SWHwAJKau56
4XJjZOiTipfRChYFr3RI6xEW8o1VqcMf0BXCC7k/Zu+yGAlCHCVDMhTJU+oMcwBX
8D3AWGQv08LBw3UrmuQF+J96M/J0v1X6Y4qcpyHmKke11nGcRorwCReWXH65NRcv
Tj3BU6ZL5ATWCx2bPBlizvKyxbHbXW4KAz5nINS7qH1cj4LIdh2nF22v759U8DT8
X8F+MeJpAH8RX9rx9Fbq1TKfB31QPLm9p4pNsVINEhBmbyccWJj8gckWIkZxVDvg
IujJ/+eMo/AkMKQcD8O/AimKcw+HV0+iRcSrPZnj0HU6p3dmKllqVHIJabg5UQNB
DIunoxujjI67StjhHEvnffBTE6Jd/KZ8N/ZZX9p5aV+vLG09sJtnb5zgqUQd5ukg
yH73a6nhd5VrrF+A4whaiJ/gjDDSNgEfXlk3AA5pRU2vnUtiO02rjpIA6v1HUUGR
5dMaHlnVx0XHstFQ1jV6ehepw2cuDXn8/rRLi/yCjgeOV6Dk5ygxUGtytCJJzK0e
Tl1xSc3vkFSWz7ahUrF4Ze+x9MHFFX2/0U6JOvyvJY1mWBzvkpck6cnfWQqJascY
g9f5pFjdNkBY03phipJirOquclRSRtzbryBxsJi2WO+GPIuB+Cu2PUsKl7m8lIZd
iYcHlrQxcKFoShXhOU4wMJq0GC1Xe3jXJP8KC4oyWjcZI6XPkcJZUhsGv8FCeMWd
EtJI9efX3H1FbCIe4Q3JevtiYIzFlDH/RenTVBdDjWxLajRRlMT5vl6yY4EviCRN
TvNbH7tQYY4wfc3bCtuvC5CgaI9u8xLAkZchvfj1XUVb5HCz7zkZ8oCykuaUMPkc
fF77uB2L2KPDfqynlXcbZSqIOX/EhDmDh7B/o3Wlm0ySBUbBTB1BCqfOOAOfFqpP
fkM8EPhVWPSRU7SQNFYMe9XQlDPTSLf70XTERzhYVCIE1X4k0gj4SXA2eCzSsNSH
X3lh+hAECP1OLXefGVKpSq6qtdgGlmoNab0coWzGrBATpUKtVdJm5r/gAKCjYwcR
Zx+ov7sAvKatRIfUBBo4Jy/go6zMeKXXDptXhFHb+RLb2aSlwY3VPRVnEWlAIwzJ
LaH4LLsSisoSXpEgwwgRWSKSivp34AV1ysw+ayx9vwvU2MjNI2GQ3ZNqgy7gkdUs
dFR8elbm24Ozdx4dmoke+ExFe6mfYJUNnLRaFxP2hxyjQhLfz5CGCAZ8/XC93GYx
6Vp3Z7uzn/9OOscuI96G2YITu6KGZHnHflx4qRXkFxYAIwxeglN+TqOIVJjRf02+
IoJuhHXOgQV0XvyTQa10nmuoJVj5j3O2guVFjsL1peaWhnVYOCmYMMRmgJFqULt+
g0fKROtOSuAkAjG2q2b23lu1Pk55/Smfo+bQmVC7i/RUF3+VbE045Nhwp3iZd+do
qdtwi8rg2yQaFK85KpgCm4TWFknDY853qXgZddrKUPJmMgAFegoOtGwVqt3iApf0
0nCFea4w9REwHi2YSOe8/Gkz5OoLqKeche0B/A8He7oTqOaFwzEPM2JSh2jn46jw
fajBaLdUDV+yO8PG/CVCBJxR8mqfnhxWv4rzrloLid08HygWgPwXp4Sz7nTWWenN
/ju7+iHfSHoLRRXsBQXMDRsAEsPQaCarBKx0DGNbbRB1cJVa5C34AE6022sNKgqw
Ym7naSh4GeLqVNM4rJvs9hrRPyKv2Gx18Gh8/LdTggGiV22QtCzj0dmD1Gh5tE/1
FKJYsWSBMkA96v9yMygOMUwbR0r+qkKLOQ/jMeM5VRBSAJCm57D1Lc4RnGZUzE7Z
8AVqeIDwS4n1SruRZkRphflpTRZ14WfBrs7ol3mzUuB0tvLTySA1T1KjMmtZlJk0
7ZhuMWONaiEGP7J2pdhrZgB3ypUffbWpnicyL4lI8RuGONlo1thjTHxiWIp/o2Gc
pCnbMET/LV+uDjJ4j1pqPvVYLQmRFe6tWJ3O2MB4O8wly8xVeNh2mjQ+gbXbnvLm
kLOVQL6vZSCnM1ouckSCr3X/AjGoYVztkG074ycyTHmJdIq+cE81J8yRYC5aGUH0
Z0sCGlCXe5q0tV7z2TjEHeVk3EXH+0PCXt81AZtT8S6mpl2kXFrFhVP4DAFKi1F/
IgfA6Cc05enxKY8XsV1d3l4QrPN9KnSCtilThKG4ZBHghWAHyBJu+VgTsciWWUBC
Le46qxW48y9NhAqOKVYZeiswxVeTZ5kejchvKhj+tt42LsISwXztMTwj/ybs1hNE
AQ4Yj2Pur3hy9FXhoiyWj+JBtJH9r1TpiKgB/Jtmm+t/ulL+gfGWeK5/B//EqHN+
oV8VLomv3QDiagrUsDLtC7J9RDzsme2zgDjOVDrHlYFy8J4D04uDn11g+Gx/tjnW
qeOR6YDlIYr/+Bt9atc2VpG8AETFqKUW73+S4MrLFq/Sjb1AqiKVBWPM8R7aYi7e
fFgaJ+d+8z3BrK7ATgn3CGRKke9Rw4/B9kBzus66r2pnga/fInHBizCjacVUo03w
UpZpjL3CifWlTec4Mo+8Hh2UN1AhAnxtF5vOoQNnaV1nTv1w3gvsa+tzNvzYCuCr
Nzrur1ashu+xpaBI2xYPW+1CDa94GUoUXJAk2nRvpA0tH//xR2Iik+nKTQTAaZCn
B34sJhc0J1W8QikVmkWhhdcdTibpoBhPiqX6mH1cJlA2HAZQHxGLRZlbq6bHcdAK
AuFZTU5jOEM/grj0QcJX8gLO/Ehs+5ew7mliY2YoDyPBz/RMUwaUbK3AP+O3NSTf
CK6prOVOL7g2RyMOtDKFfH7LuYDbAf9oDMkk9XvcBWlZssQNP0XH6vI1JsI/XLoM
enJp6mM7xvxIUDCG+WYmfru5SxX3iN3uVvyEv64xqBWiCkMP9lmGli+0ci8yjLqO
rjZ1mzaeR12DZ4oFHFR5nWF1f12m51uXQqw0BxgC0IAoOB/C6IcTGWWHa5A2N338
FlM0W43HF6vEQkPFrvFHcl4brlv3qYsLE0fQnvM9LN6WP3A8Oe+dBNQSuu9Urk4N
ncXw0sDAGWqV6yy5RzAHbtVO5jAmarZS0QuPK0mOQkf6QIDQkOGpy6BIs3enksTb
ttpW0ajTc4Vnl+rEDs1+8e2zR5Uhfn4X1HhdQ748sUvlfxnlWnTUyPaF3knc5PmR
qccyVokd4/dZGMh3kbJbW+wdpcARwZSidNSivknU39flep2WG5+zS7FwCSV9sXH6
P7nfHvPj39uYONVDoERdzzcbt4a1GbJ/T1eT6rI1f22zU3d0fNSNF9a5JjjaVy5P
WLc4tnVGXdgxfylGZj5oRtCz6/ZzQk3QqVE+Qj9G7IEXXHYQZ4TVzHw/vmUZErck
ngE28zmGk66opDPh5TOX7AKD7ZU8lfqqQod2QD+7fw3BrsXj+h5EKhNBsL28QufL
eMaz9cnGE69uN8S9e4HNjbHFiTteJ1xWNdz5VYuEL5LobNhrQiMLPUBjaOuQvNLp
M+v/MqiHaYKHY0pFZHkiYy1dy9wg3S2WcdO5tWbvnGvHuIMFuq3K+38otAJuc9W5
0UnBiNk3hYpcwjhphHd4z+wIO3vIaHSg09gOc5APlmd8INRzUZNGz0PB8gvoKl56
US0vs9cozTFfR73+gpcGaVepOhnEtZw50d702FUCrMTjNiYv/DrRMCPhpuQRnfwC
jq3JqPGvAL1+IUsNsSBZMo0KQ7G+Xy7vlOiboPrvBctAsPOxE8bNFnUw2moCbvXk
3dUa0FNerwgSufLNEECgyqH9MBmiW3FbgfH6GwR0E84QHbGSzyaA4EBt6RmUJFPq
m5JdwlQeqy5zcC7iBD81qlwNsRjTH/5934Xc4wgmaaYrxxj0oGfB5yTr2IGDmKnU
dIjzMAMnr5PubrpXPfDuIvlpbSflyNJczp7m4dkzlr6iT95bOT+oXKfPkLzGDVqG
dcHHHYna3YEmMGNvOW3uHuswIMbUiiziLiTym5/RryCNbRdMk+A9q6HfVlQi6Eg0
HjsnTKtd/iTE7JKebsTQJ73x+LCaeidWmpojUyjWE76tU3y36jLy1N5P+07qr6Q3
NhnJs2SKC1aVU1720sztPZ6yoh8S/AE8pC8+Gu5Un08AyXlysE/Zo/bCILiGBBN3
KraROOYdj5DiJlgl9Ut2uNhfIQpK02vbFHN0E7++62+gQ15o0a4vy940dK7NNsaL
yHAcN+wF1issJgMrqEGwWRoW3ROmEf7S3hZc5W7G009wlO3cmISIgoRwAEaS0SG6
U3H25DP4exdRq2qEHUqvAOeUPNz2MnO9+0eaFpyhbTf5NAw3Bp5lzu3YL21m0OIL
+OAUfTpZcmFCAKeO8BeGgcF6sNUeMjoY1SVxjTkA/zb9dy9a6ZM6bFI8zykgO81N
T1jIPDFqHz8Xjy5+kKViZ81Y8unjWlkS8RuhrsYKzguXAQfMoDZDoTzaMaDmCPNB
/8EzaLZPLvef2GXe4u+KXGoI6dbicCZSFpBvgG6YVDQrRXKbqQbOGRXibAVnNPBf
mG1WUBIArMLPgjOlGFS2OACEmf7zB/yRn9MAB9HgEpjSXm28YcVpYp3ypQ17STaD
CL5Yanh0HCWLNTqJEWhopE+xp3AQgFao7OVdileGnw3KX4AQdl0ERQJfNwFEEPMX
4vMC6dSmKLKdER+i3CPSQFniLbqkyPvJJSgkHyD7wXg/RLP9g27iS9hbwIF5rNlW
y7jLJE3sWzvtYR9wosUaG0g62qcsbwiX3UtQSag2Cx1MDnoh8nz5vzf3SAy42tZt
3tXsN12WyhwsloU2sSWfBgX1dopl1C8E01/kqydJensb3jXhxYFcZ+mc8C1AX2Q9
ItP+wCft4IMrPHS9zYPttyCedF8MKBwcFhBN5N5AN0ypxdz4W7vE+mGTnrKEiuwE
7tTQHybJnVByg3pIz03sl7QExBvkG4cQfGZPNQumQj26cZ1FjZvBsTjgEDypGfFB
bxdjShhn0byZdf1AFSTVvcYdtlZZIQsCYbQFhH3zObwXhZKDbl2MUbWcT+NqBzk5
5inTBpc1XdJrMgsN0oAkSajp5STSkVseTmZzWen0eEEWm1IRwJMzO01sfMjde2uq
sEtorSWodfY/RcNuu6WE5qUs0eSlCD+HpwnO8ueQAKJcguzqx5pM/uvQ+nqIKQ8U
Eaf4ama45Eacd4ZUpHRJ2GGdQL3kk1qAUmUbvJMjW+jhNiCANJEv3Tj2C5P7cxMJ
ghbzWKeDJkKT8n7vhFjbRPpE7FZz8iFvwGXV0VwJ11TeDrEIslbhPcqKlDxA0imY
jI+TKkIBfHe4hU11mv0+7Z1f/OpVACd8AQOzhUW3IvsLWGbAMryPte6LgtHCFLuV
h/5+qjQ0Kf8G/ON/4LEzB5nd4xCJCXqR1DOjUgctsFpwPOz387TunIy9oG4XCJqb
+Ddbm94JcTuAthH7F5Yo/p4DmsnXCKZJS60B7MEOnzg2ohA225d1GeW09IvO0icc
13unBrVIPVsrn073ceFZLeaZEJXMmppNvgVaOJTuELCv7vuCW8gOwAWXTNVFDIl+
GTLQGgwX/WyNujjIMNDQa+rpFcHd26/ltpvKbMqKRz3Nw29dMUle3AqoXl9UMSs3
yDq0K3z2xumOqPKNf06HPu1S+fk1o92AdoJsiG7KpDtZUHtwf2iVO87kQxHJ7wz5
ntwrRjeUlSyjeed+vwTWPCIVopVgdvfJl+ZAPRNXYJC3ilkPQzsJoc0VRUTM6Hk5
EN+HBFrqMSe3dFDY5U/nmnlHRD5U6l+OYxx/PkHzwnmcwZTCHaOykTNmwbqTKwdb
VPmfjKjj+17wmUCf85uj0G/UWxytokQmWPmrK5N5r/6VQfXObOMyCZ/RJVzNkc4m
3UTednJCO3qCoHbwpOszEdRdxIkPniEQCMgmEk80yeXW+8k68HFvF0GwwjENM9Mu
4PayrVDXj0+Z5NP4CMNOXU3Qk97ZsmG5SWB+5TrqnwJknRkIkLhbn+VJEj8BFEYP
qchXylh8ve4BDrWz/fcbYOrAG2noQcJ4DYNJWEZJQiMZEhJXUY0ERQmUdA/pwcm0
P3ZeUTXPgylFEDnmVphnULQUO8hIHPHVVuBcydFj9P70850gvw6QnsBPg/BVzHpH
jMAp90JvhI/kc0Ws8sbtUMpcBEPWNx7NZ3/TUL3ZX/MHOpKYtAEdLG//yk1iLiBD
`pragma protect end_protected
