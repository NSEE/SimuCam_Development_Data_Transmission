package avalon_mm_data_buffer_pkg is
	
end package avalon_mm_data_buffer_pkg;

package body avalon_mm_data_buffer_pkg is
	
end package body avalon_mm_data_buffer_pkg;
