library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity data_controller_ent is
	port(
		clk : in std_logic;
		rst : in std_logic
	);
end entity data_controller_ent;

architecture RTL of data_controller_ent is
	
begin

end architecture RTL;
